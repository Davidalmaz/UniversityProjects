CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 1 100 9
1 79 585 671
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
16 C:\CM60S\BOM.DAT
0 7
1 79 585 671
143654930 0
0
6 Title:
5 Name:
0
0
0
18
13 Logic Switch~
5 172 294 0 1 11
0 7
0
0 0 21360 0
2 0V
-6 -16 8 -8
1 D
-3 -26 4 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
8953 0 0
0
0
13 Logic Switch~
5 172 334 0 1 11
0 6
0
0 0 21360 0
2 0V
-6 -16 8 -8
1 C
-3 -26 4 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
4441 0 0
0
0
13 Logic Switch~
5 173 372 0 1 11
0 5
0
0 0 21360 0
2 0V
-6 -16 8 -8
1 B
-3 -26 4 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3618 0 0
0
0
13 Logic Switch~
5 172 414 0 1 11
0 4
0
0 0 21360 0
2 0V
-6 -16 8 -8
1 A
-3 -26 4 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
6153 0 0
0
0
13 Logic Switch~
5 159 180 0 10 11
0 8 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
7 Despeje
-23 -26 26 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
5394 0 0
0
0
13 Logic Switch~
5 225 157 0 10 11
0 3 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
5 Carga
-16 -26 19 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
7734 0 0
0
0
13 Logic Switch~
5 224 211 0 10 11
0 12 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
6 Conteo
-20 -26 22 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
9914 0 0
0
0
7 Pulser~
4 114 268 0 10 12
0 15 16 9 17 0 0 5 5 3
7
0
0 0 4656 0
0
3 CLK
-10 -28 11 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
1 V
3747 0 0
0
0
10 2-In NAND~
219 395 389 0 3 22
0 10 11 18
0
0 0 624 180
6 74LS00
-14 -24 28 -16
3 U2A
-8 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 512 4 1 1 0
1 U
3549 0 0
0
0
7 74LS161
96 301 278 0 14 29
0 12 12 9 7 6 5 4 3 8
19 11 13 10 14
0
0 0 13040 0
8 74LS161A
-28 -60 28 -52
2 U1
-7 -61 7 -53
0
15 DVCC=16;DGND=8;
126 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 7 10 2 6 5 4 3 9 1
15 11 12 13 14 7 10 2 6 5
4 3 9 1 15 11 12 13 14 0
65 0 0 512 1 0 0 0
1 U
7931 0 0
0
0
7 Ground~
168 473 87 0 1 3
0 2
0
0 0 53360 0
0
4 GND4
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
9325 0 0
0
0
7 Ground~
168 423 87 0 1 3
0 2
0
0 0 53360 0
0
4 GND3
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
8903 0 0
0
0
7 Ground~
168 363 90 0 1 3
0 2
0
0 0 53360 0
0
4 GND2
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3834 0 0
0
0
7 Ground~
168 306 89 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3363 0 0
0
0
5 Lamp~
206 463 68 0 2 3
11 14 2
0
0 0 608 0
3 100
-10 -24 11 -16
1 A
-4 -22 3 -14
0
0
11 %D %1 %2 %V
0
0
0
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 L
7668 0 0
0
0
5 Lamp~
206 410 68 0 2 3
11 10 2
0
0 0 608 0
3 100
-10 -24 11 -16
1 B
-4 -22 3 -14
0
0
11 %D %1 %2 %V
0
0
0
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 L
4718 0 0
0
0
5 Lamp~
206 351 70 0 2 3
11 13 2
0
0 0 608 0
3 100
-10 -24 11 -16
1 C
-4 -22 3 -14
0
0
11 %D %1 %2 %V
0
0
0
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 L
3874 0 0
0
0
5 Lamp~
206 295 70 0 2 3
11 11 2
0
0 0 608 0
3 100
-10 -24 11 -16
1 D
-4 -22 3 -14
0
0
11 %D %1 %2 %V
0
0
0
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 L
6671 0 0
0
0
19
1 8 3 0 0 4224 0 6 10 0 0 4
237 157
343 157
343 242
339 242
1 7 4 0 0 8320 0 4 10 0 0 4
184 414
229 414
229 314
269 314
1 6 5 0 0 8320 0 3 10 0 0 4
185 372
216 372
216 305
269 305
1 5 6 0 0 12416 0 2 10 0 0 4
184 334
205 334
205 296
269 296
1 4 7 0 0 8320 0 1 10 0 0 3
184 294
184 287
269 287
9 1 8 0 0 12432 0 10 5 0 0 4
339 251
353 251
353 180
171 180
3 3 9 0 0 8320 0 10 8 0 0 3
269 260
269 259
138 259
0 1 10 0 0 8192 0 0 9 14 0 4
393 305
472 305
472 398
419 398
0 2 11 0 0 8192 0 0 9 12 0 5
355 287
355 341
429 341
429 380
419 380
2 0 12 0 0 8192 0 10 0 0 11 3
269 251
261 251
261 242
1 1 12 0 0 8320 0 7 10 0 0 4
236 211
261 211
261 242
269 242
1 11 11 0 0 16512 0 18 10 0 0 6
283 83
275 83
275 124
362 124
362 287
333 287
12 1 13 0 0 8320 0 10 17 0 0 5
333 296
377 296
377 112
339 112
339 83
13 1 10 0 0 8320 0 10 16 0 0 4
333 305
393 305
393 81
398 81
14 1 14 0 0 8320 0 10 15 0 0 5
333 314
405 314
405 110
451 110
451 81
1 2 2 0 0 4224 0 11 15 0 0 2
473 81
475 81
1 2 2 0 0 0 0 12 16 0 0 2
423 81
422 81
1 2 2 0 0 0 0 13 17 0 0 2
363 84
363 83
1 2 2 0 0 0 0 14 18 0 0 2
306 83
307 83
0
0
2049 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
592328 1210432 100 100 0 0
0 0 0 0
2 74 163 144
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
12385 0
4 1 2
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
