CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 9
32 88 1248 655
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
16 C:\CM60S\BOM.DAT
0 7
32 88 1248 655
143654930 0
0
6 Title:
5 Name:
0
0
0
18
13 Logic Switch~
5 147 281 0 10 11
0 10 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
1 D
-3 -26 4 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
8953 0 0
0
0
13 Logic Switch~
5 150 217 0 1 11
0 11
0
0 0 21360 0
2 0V
-6 -16 8 -8
1 C
-3 -26 4 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
4441 0 0
0
0
13 Logic Switch~
5 146 146 0 10 11
0 12 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
1 B
-3 -26 4 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3618 0 0
0
0
13 Logic Switch~
5 145 83 0 10 11
0 9 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-5 -15 9 -7
1 A
-3 -26 4 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
6153 0 0
0
0
7 Ground~
168 520 359 0 1 3
0 2
0
0 0 53360 0
0
4 GND2
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
5394 0 0
0
0
10 3-In NAND~
219 470 354 0 4 22
0 6 5 4 3
0
0 0 624 0
6 74LS10
-21 -28 21 -20
3 U2C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
17

0 9 10 11 8 1 2 13 12 3
4 5 6 9 10 11 8 0
65 0 0 0 3 3 2 0
1 U
7734 0 0
0
0
10 3-In NAND~
219 380 297 0 4 22
0 9 8 7 6
0
0 0 624 0
6 74LS10
-21 -28 21 -20
3 U2B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
17

0 3 4 5 6 1 2 13 12 3
4 5 6 9 10 11 8 0
65 0 0 0 3 2 2 0
1 U
9914 0 0
0
0
10 2-In NAND~
219 300 405 0 3 22
0 11 10 4
0
0 0 624 0
6 74LS00
-14 -24 28 -16
3 U3C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 3 0
1 U
3747 0 0
0
0
10 2-In NAND~
219 301 346 0 3 22
0 12 10 5
0
0 0 624 0
6 74LS00
-14 -24 28 -16
3 U3B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 3 0
1 U
3549 0 0
0
0
7 Ground~
168 478 170 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
7931 0 0
0
0
10 2-In NAND~
219 231 284 0 3 22
0 10 10 7
0
0 0 624 0
6 74LS00
-14 -24 28 -16
3 U3A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 3 0
1 U
9325 0 0
0
0
10 2-In NAND~
219 233 135 0 3 22
0 12 12 8
0
0 0 624 0
6 74LS00
-14 -24 28 -16
3 U1D
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 1 0
1 U
8903 0 0
0
0
10 2-In NAND~
219 435 164 0 3 22
0 14 15 13
0
0 0 624 0
6 74LS00
-14 -24 28 -16
3 U1C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 1 0
1 U
3834 0 0
0
0
10 3-In NAND~
219 310 93 0 4 22
0 9 8 7 14
0
0 0 624 0
6 74LS10
-21 -28 21 -20
3 U2A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
17

0 1 2 13 12 1 2 13 12 3
4 5 6 9 10 11 8 0
65 0 0 0 3 1 2 0
1 U
3363 0 0
0
0
10 2-In NAND~
219 344 235 0 3 22
0 16 16 15
0
0 0 624 0
6 74LS00
-14 -24 28 -16
3 U1B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 1 0
1 U
7668 0 0
0
0
10 2-In NAND~
219 240 226 0 3 22
0 11 11 16
0
0 0 624 0
6 74LS00
-14 -24 28 -16
3 U1A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 1 0
1 U
4718 0 0
0
0
5 Lamp~
206 510 340 0 2 3
11 3 2
0
0 0 624 0
3 100
-10 -24 11 -16
2 L2
-7 -22 7 -14
0
0
11 %D %1 %2 %V
0
0
0
5

0 1 2 1 2 0
82 0 0 0 0 0 0 0
1 L
3874 0 0
0
0
5 Lamp~
206 468 151 0 2 3
11 13 2
0
0 0 624 0
3 100
-10 -24 11 -16
2 L1
-7 -22 7 -14
0
0
11 %D %1 %2 %V
0
0
0
5

0 1 2 1 2 0
82 0 0 0 0 0 0 0
1 L
6671 0 0
0
0
28
4 0 3 0 0 4096 0 6 0 0 3 2
497 354
498 353
1 2 2 0 0 4240 0 5 17 0 0 2
520 353
522 353
1 3 3 0 0 4240 0 17 0 0 0 2
498 353
504 353
3 3 4 0 0 4224 0 6 8 0 0 4
446 363
335 363
335 405
327 405
2 3 5 0 0 4224 0 6 9 0 0 4
446 354
336 354
336 346
328 346
4 1 6 0 0 8320 0 7 6 0 0 4
407 297
438 297
438 345
446 345
0 3 7 0 0 8192 0 0 7 16 0 3
278 284
278 306
356 306
0 2 8 0 0 4224 0 0 7 17 0 3
270 135
270 297
356 297
0 1 9 0 0 12416 0 0 7 24 0 5
262 83
262 116
291 116
291 288
356 288
0 2 10 0 0 4224 0 0 8 21 0 3
181 281
181 414
276 414
0 1 11 0 0 4224 0 0 8 28 0 3
191 217
191 396
276 396
0 2 10 0 0 0 0 0 9 21 0 3
186 281
186 355
277 355
0 1 12 0 0 4224 0 0 9 19 0 3
175 146
175 337
277 337
1 2 2 0 0 128 0 10 18 0 0 2
478 164
480 164
1 3 13 0 0 4224 0 18 13 0 0 2
456 164
462 164
3 3 7 0 0 8320 0 11 14 0 0 4
258 284
278 284
278 102
286 102
3 2 8 0 0 128 0 12 14 0 0 4
260 135
278 135
278 93
286 93
2 0 12 0 0 0 0 12 0 0 19 3
209 144
209 146
201 146
1 1 12 0 0 128 0 3 12 0 0 4
158 146
201 146
201 126
209 126
2 0 10 0 0 0 0 11 0 0 21 3
207 293
196 293
196 281
1 1 10 0 0 128 0 1 11 0 0 4
159 281
199 281
199 275
207 275
4 1 14 0 0 4224 0 14 13 0 0 4
337 93
403 93
403 155
411 155
3 2 15 0 0 8320 0 15 13 0 0 4
371 235
403 235
403 173
411 173
1 1 9 0 0 128 0 4 14 0 0 4
157 83
279 83
279 84
286 84
2 0 16 0 0 8192 0 15 0 0 27 3
320 244
308 244
308 226
2 0 11 0 0 0 0 16 0 0 28 3
216 235
204 235
204 217
1 3 16 0 0 4224 0 15 16 0 0 2
320 226
267 226
1 1 11 0 0 128 0 2 16 0 0 2
162 217
216 217
0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
