CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 70 30 100 9
4 82 836 649
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
16 C:\CM60S\BOM.DAT
0 7
4 82 836 649
143654930 0
0
6 Title:
5 Name:
0
0
0
24
13 Logic Switch~
5 223 303 0 10 11
0 15 0 0 0 0 0 0 0 0
1
0
0 0 21344 0
2 5V
-6 -16 8 -8
1 D
-3 -26 4 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
8953 0 0
0
0
13 Logic Switch~
5 226 244 0 1 11
0 13
0
0 0 21344 0
2 0V
-6 -16 8 -8
1 C
-3 -26 4 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
4441 0 0
0
0
13 Logic Switch~
5 227 184 0 1 11
0 5
0
0 0 21344 0
2 0V
-6 -16 8 -8
1 B
-3 -26 4 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
3618 0 0
0
0
13 Logic Switch~
5 226 116 0 10 11
0 6 0 0 0 0 0 0 0 0
1
0
0 0 21344 0
2 5V
-6 -16 8 -8
1 A
-3 -26 4 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
6153 0 0
0
0
10 2-In NAND~
219 416 409 0 3 22
0 4 3 12
0
0 0 608 0
6 74LS00
-14 -24 28 -16
3 U4C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 4 0
1 U
5394 0 0
0
0
10 2-In NAND~
219 327 435 0 3 22
0 6 13 3
0
0 0 608 0
6 74LS00
-14 -24 28 -16
3 U4B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 4 0
1 U
7734 0 0
0
0
10 2-In NAND~
219 324 372 0 3 22
0 6 5 4
0
0 0 608 0
6 74LS00
-14 -24 28 -16
3 U4A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 4 0
1 U
9914 0 0
0
0
7 Ground~
168 514 270 0 1 3
0 2
0
0 0 53344 0
0
4 GND3
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3747 0 0
0
0
9 Inverter~
13 464 138 0 2 22
0 7 8
0
0 0 608 0
6 74LS04
-21 -19 21 -11
3 U1E
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 11 10 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 5 1 0
1 U
3549 0 0
0
0
10 3-In NAND~
219 415 177 0 4 22
0 11 10 9 7
0
0 0 608 0
6 74LS10
-21 -28 21 -20
3 U2A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
17

0 1 2 13 12 1 2 13 12 3
4 5 6 9 10 11 8 0
65 0 0 0 3 1 2 0
1 U
7931 0 0
0
0
7 Ground~
168 697 258 0 1 3
0 2
0
0 0 53344 0
0
4 GND5
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
9325 0 0
0
0
7 Ground~
168 502 336 0 1 3
0 2
0
0 0 53344 0
0
4 GND4
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
8903 0 0
0
0
7 Ground~
168 527 198 0 1 3
0 2
0
0 0 53344 0
0
4 GND2
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3834 0 0
0
0
7 Ground~
168 504 117 0 1 3
0 2
0
0 0 53344 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3363 0 0
0
0
9 2-In XOR~
219 412 252 0 3 22
0 5 13 16
0
0 0 608 0
6 74LS86
-21 -24 21 -16
3 U3A
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 3 0
1 U
7668 0 0
0
0
9 Inverter~
13 324 317 0 2 22
0 15 14
0
0 0 608 0
6 74LS04
-21 -19 21 -11
3 U1D
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 9 8 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 4 1 0
1 U
4718 0 0
0
0
9 Inverter~
13 326 253 0 2 22
0 13 9
0
0 0 608 0
6 74LS04
-21 -19 21 -11
3 U1C
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 1 0
1 U
3874 0 0
0
0
9 Inverter~
13 327 189 0 2 22
0 5 10
0
0 0 608 0
6 74LS04
-21 -19 21 -11
3 U1B
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 1 0
1 U
6671 0 0
0
0
9 Inverter~
13 333 129 0 2 22
0 6 11
0
0 0 608 0
6 74LS04
-21 -19 21 -11
3 U1A
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 1 0
1 U
3789 0 0
0
0
5 Lamp~
206 687 239 0 2 3
11 12 2
0
0 0 624 0
3 100
-10 -24 11 -16
2 L5
-7 -22 7 -14
0
0
11 %D %1 %2 %V
0
0
0
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 L
4871 0 0
0
0
5 Lamp~
206 492 317 0 2 3
11 14 2
0
0 0 624 0
3 100
-10 -24 11 -16
2 L4
-7 -22 7 -14
0
0
11 %D %1 %2 %V
0
0
0
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 L
3750 0 0
0
0
5 Lamp~
206 503 251 0 2 3
11 13 2
0
0 0 624 0
3 100
-10 -24 11 -16
2 L3
-7 -22 7 -14
0
0
11 %D %1 %2 %V
0
0
0
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 L
8778 0 0
0
0
5 Lamp~
206 508 173 0 2 3
11 16 2
0
0 0 624 0
3 100
-10 -24 11 -16
2 L2
-7 -22 7 -14
0
0
11 %D %1 %2 %V
0
0
0
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 L
538 0 0
0
0
5 Lamp~
206 492 98 0 2 3
11 8 2
0
0 0 624 0
3 100
-10 -24 11 -16
2 L1
-7 -22 7 -14
0
0
11 %D %1 %2 %V
0
0
0
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 L
6843 0 0
0
0
34
2 0 3 0 0 0 0 5 0 0 14 2
392 418
392 418
1 0 4 0 0 0 0 5 0 0 13 2
392 400
392 400
3 0 3 0 0 4096 0 6 0 0 14 2
354 435
354 436
2 0 5 0 0 4096 0 7 0 0 17 2
300 381
300 382
1 0 6 0 0 4096 0 7 0 0 18 2
300 363
300 364
4 1 7 0 0 8320 0 10 9 0 0 4
442 177
446 177
446 138
449 138
1 2 2 0 0 4096 0 8 22 0 0 2
514 264
515 264
2 1 8 0 0 4224 0 9 24 0 0 3
485 138
485 111
480 111
3 0 9 0 0 0 0 10 0 0 31 2
391 186
391 186
2 0 10 0 0 0 0 10 0 0 30 2
391 177
391 177
1 0 11 0 0 0 0 10 0 0 29 2
391 168
391 168
3 1 12 0 0 4224 0 5 20 0 0 4
443 409
667 409
667 252
675 252
3 0 4 0 0 8320 0 7 0 0 0 5
351 372
351 373
388 373
388 400
396 400
0 0 3 0 0 8320 0 0 0 0 0 5
351 435
351 436
388 436
388 418
396 418
0 2 13 0 0 4224 0 0 6 32 0 5
253 244
253 445
306 445
306 444
303 444
0 1 6 0 0 4096 0 0 6 18 0 5
292 364
292 427
306 427
306 426
303 426
0 0 5 0 0 4240 0 0 0 33 0 3
267 184
267 382
305 382
0 0 6 0 0 4224 0 0 0 34 0 3
259 116
259 364
305 364
1 2 2 0 0 4096 0 11 20 0 0 2
697 252
699 252
1 2 2 0 0 0 0 12 21 0 0 2
502 330
504 330
1 2 2 0 0 8320 0 13 23 0 0 3
527 192
527 186
520 186
1 2 2 0 0 0 0 14 24 0 0 2
504 111
504 111
2 1 14 0 0 4224 0 16 21 0 0 4
345 317
472 317
472 330
480 330
1 1 15 0 0 4224 0 1 16 0 0 4
235 303
301 303
301 317
309 317
0 1 13 0 0 0 0 0 22 27 0 5
371 268
371 278
474 278
474 264
491 264
3 1 16 0 0 8320 0 15 23 0 0 4
445 252
470 252
470 186
496 186
0 2 13 0 0 0 0 0 15 32 0 3
279 244
279 261
396 261
0 1 5 0 0 0 0 0 15 33 0 5
282 184
282 213
375 213
375 243
396 243
2 0 11 0 0 8320 0 19 0 0 0 4
354 129
387 129
387 168
395 168
2 0 10 0 0 8320 0 18 0 0 0 3
348 189
348 177
395 177
2 0 9 0 0 8320 0 17 0 0 0 4
347 253
387 253
387 186
395 186
1 1 13 0 0 0 0 2 17 0 0 4
238 244
303 244
303 253
311 253
1 1 5 0 0 0 0 3 18 0 0 4
239 184
304 184
304 189
312 189
1 1 6 0 0 0 0 4 19 0 0 4
238 116
310 116
310 129
318 129
0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
