CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 5 100 9
7 86 715 789
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
16 C:\CM60S\BOM.DAT
0 7
8 362 681 505
160432146 0
0
6 Title:
5 Name:
0
0
0
8
9 2-In AND~
219 486 116 0 3 22
0 6 3 5
0
0 0 608 0
6 74LS08
-21 -24 21 -16
3 AND
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 1 0
1 U
8953 0 0
0
0
5 SCOPE
12 545 105 0 1 11
0 5
0
0 0 57568 0
3 SAL
-11 -4 10 4
2 U2
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
0
4441 0 0
0
0
5 SCOPE
12 389 132 0 1 11
0 3
0
0 0 57568 0
2 E1
-7 -4 7 4
2 U2
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
0
3618 0 0
0
0
5 SCOPE
12 389 106 0 1 11
0 6
0
0 0 57568 0
2 E2
-8 -4 6 4
2 U2
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
0
6153 0 0
0
0
7 Ground~
168 362 192 0 1 3
0 2
0
0 0 53344 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
5394 0 0
0
0
7 Pulser~
4 125 126 0 10 12
0 7 8 4 9 0 0 5 5 3
7
0
0 0 4640 0
0
5 RELOJ
-17 -28 18 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
1 V
7734 0 0
0
0
6 74LS93
109 281 108 0 8 17
0 2 2 4 3 10 11 6 3
0
0 0 13024 0
6 74LS93
-21 -35 21 -27
4 CONT
-14 -36 14 -28
0
15 DVCC=5;DGND=10;
76 %D [%5bi %10bi %1i %2i %3i %4i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o] %M
0
12 type:digital
5 DIP14
17

0 2 3 14 1 11 8 9 12 2
3 14 1 11 8 9 12 0
65 0 0 512 1 0 0 0
1 U
9914 0 0
0
0
5 Lamp~
206 595 103 0 2 3
11 5 2
0
0 0 608 0
3 100
-10 -24 11 -16
4 LAMP
-14 -22 14 -14
0
0
11 %D %1 %2 %V
0
0
0
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 L
3747 0 0
0
0
11
2 1 2 0 0 12416 0 8 5 0 0 5
607 116
611 116
611 178
362 178
362 186
4 8 3 0 0 12288 0 7 7 0 0 5
243 126
239 126
239 155
313 155
313 126
3 3 4 0 0 4224 0 6 7 0 0 2
149 117
243 117
1 0 5 0 0 4096 0 2 0 0 11 2
545 117
545 116
1 0 3 0 0 0 0 3 0 0 8 2
389 144
389 145
1 0 6 0 0 4096 0 4 0 0 7 2
389 118
389 117
7 1 6 0 0 4224 0 7 1 0 0 6
313 117
456 117
456 107
463 107
463 107
462 107
8 2 3 0 0 12416 0 7 1 0 0 8
313 126
325 126
325 145
456 145
456 125
463 125
463 125
462 125
2 0 2 0 0 0 0 7 0 0 10 2
249 108
225 108
1 1 2 0 0 0 0 7 5 0 0 5
249 99
225 99
225 178
362 178
362 186
3 1 5 0 0 4224 0 1 8 0 0 2
507 116
583 116
0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
