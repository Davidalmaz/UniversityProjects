CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 9
0 71 1280 672
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
16 C:\CM60S\BOM.DAT
0 7
0 71 1280 672
143654930 0
0
6 Title:
5 Name:
0
0
0
18
13 Logic Switch~
5 215 374 0 10 11
0 12 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V5
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
8953 0 0
0
0
13 Logic Switch~
5 198 332 0 1 11
0 4
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V4
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
4441 0 0
0
0
13 Logic Switch~
5 196 282 0 10 11
0 5 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V3
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
3618 0 0
0
0
13 Logic Switch~
5 193 224 0 10 11
0 6 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
6153 0 0
0
0
13 Logic Switch~
5 192 167 0 10 11
0 7 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
5394 0 0
0
0
9 2-In XOR~
219 312 301 0 3 22
0 4 12 8
0
0 0 624 0
6 74LS86
-21 -24 21 -16
3 U2D
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 1 0
1 U
7734 0 0
0
0
9 2-In XOR~
219 315 259 0 3 22
0 5 12 9
0
0 0 624 0
6 74LS86
-21 -24 21 -16
3 U2C
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 1 0
1 U
9914 0 0
0
0
9 2-In XOR~
219 315 215 0 3 22
0 6 12 10
0
0 0 624 0
6 74LS86
-21 -24 21 -16
3 U2B
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 1 0
1 U
3747 0 0
0
0
9 2-In XOR~
219 317 174 0 3 22
0 7 12 11
0
0 0 624 0
6 74LS86
-21 -24 21 -16
3 U2A
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 1 0
1 U
3549 0 0
0
0
6 74LS83
105 455 149 0 14 29
0 3 2 2 3 11 10 9 8 12
17 16 15 14 13
0
0 0 13040 0
7 74LS83A
-24 -60 25 -52
2 U1
-7 -61 7 -53
0
15 DVCC=5;DGND=12;
125 %D [%5bi %12bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 3 8 10 16 4 7 11 13
15 2 6 9 14 1 3 8 10 16
4 7 11 13 15 2 6 9 14 0
65 0 0 0 1 0 0 0
1 U
7931 0 0
0
0
7 Ground~
168 659 175 0 1 3
0 2
0
0 0 53360 90
0
4 GND1
-14 -28 14 -20
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
9325 0 0
0
0
9 V Source~
197 292 100 0 2 5
0 3 2
0
0 0 17264 0
3 10V
13 0 34 8
3 Vs1
13 -10 34 -2
0
0
11 %D %1 %2 %V
0
0
0
5

0 1 2 1 2 0
86 0 0 0 1 0 0 0
2 Vs
8903 0 0
0
0
7 Ground~
168 346 130 0 1 3
0 2
0
0 0 53360 0
0
4 GND2
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3834 0 0
0
0
5 Lamp~
206 567 85 0 2 3
11 17 2
0
0 0 608 0
3 100
-10 -24 11 -16
2 s4
-7 -22 7 -14
0
0
11 %D %1 %2 %V
0
0
0
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 L
3363 0 0
0
0
5 Lamp~
206 568 125 0 2 3
11 16 2
0
0 0 608 0
3 100
-10 -24 11 -16
2 s3
-7 -22 7 -14
0
0
11 %D %1 %2 %V
0
0
0
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 L
7668 0 0
0
0
5 Lamp~
206 569 164 0 2 3
11 15 2
0
0 0 608 0
3 100
-10 -24 11 -16
2 s2
-7 -22 7 -14
0
0
11 %D %1 %2 %V
0
0
0
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 L
4718 0 0
0
0
5 Lamp~
206 569 204 0 2 3
11 14 2
0
0 0 608 0
3 100
-10 -24 11 -16
2 s1
-7 -22 7 -14
0
0
11 %D %1 %2 %V
0
0
0
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 L
3874 0 0
0
0
5 Lamp~
206 574 328 0 2 3
11 13 2
0
0 0 608 0
3 100
-10 -24 11 -16
7 ACARREO
-24 -22 25 -14
0
0
11 %D %1 %2 %V
0
0
0
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 L
6671 0 0
0
0
28
0 3 2 0 0 8192 0 0 10 2 0 3
396 122
396 131
423 131
0 2 2 0 0 8192 0 0 10 18 0 3
344 119
344 122
423 122
0 4 3 0 0 4096 0 0 10 4 0 3
383 75
383 140
423 140
1 1 3 0 0 8320 0 12 10 0 0 5
292 79
292 75
415 75
415 113
423 113
1 1 4 0 0 8320 0 2 6 0 0 5
210 332
210 291
288 291
288 292
296 292
1 1 5 0 0 8320 0 3 7 0 0 5
208 282
208 251
291 251
291 250
299 250
1 1 6 0 0 8320 0 4 8 0 0 3
205 224
205 206
299 206
1 1 7 0 0 4224 0 5 9 0 0 4
204 167
293 167
293 165
301 165
8 3 8 0 0 8320 0 10 6 0 0 4
423 176
392 176
392 301
345 301
7 3 9 0 0 8320 0 10 7 0 0 4
423 167
373 167
373 259
348 259
3 6 10 0 0 12416 0 8 10 0 0 4
348 215
362 215
362 158
423 158
3 5 11 0 0 8320 0 9 10 0 0 3
350 174
350 149
423 149
2 0 12 0 0 4096 0 6 0 0 16 2
296 310
242 310
2 0 12 0 0 4096 0 7 0 0 16 2
299 268
242 268
2 0 12 0 0 0 0 8 0 0 16 2
299 224
242 224
2 0 12 0 0 8320 0 9 0 0 17 3
301 183
242 183
242 374
1 9 12 0 0 0 0 1 10 0 0 4
227 374
415 374
415 194
423 194
2 1 2 0 0 0 0 12 13 0 0 6
292 121
292 126
333 126
333 119
346 119
346 124
2 0 2 0 0 0 0 17 0 0 21 3
581 217
620 217
620 177
2 0 2 0 0 8320 0 18 0 0 22 4
586 341
642 341
642 176
647 176
2 0 2 0 0 0 0 15 0 0 23 3
580 138
620 138
620 177
2 0 2 0 0 0 0 14 0 0 23 3
579 98
647 98
647 176
2 1 2 0 0 0 0 16 11 0 0 4
581 177
644 177
644 176
652 176
14 1 13 0 0 4224 0 10 18 0 0 3
487 194
487 341
562 341
13 1 14 0 0 8320 0 10 17 0 0 4
487 167
522 167
522 217
557 217
12 1 15 0 0 4224 0 10 16 0 0 4
487 158
549 158
549 177
557 177
11 1 16 0 0 4224 0 10 15 0 0 4
487 149
548 149
548 138
556 138
10 1 17 0 0 8320 0 10 14 0 0 3
487 140
487 98
555 98
1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 4
235 85 275 109
245 93 277 109
4 1001
0
2049 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
671286808 1079360 100 100 0 0
0 0 0 0
1 66 162 136
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
12385 0
4 1 5
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
