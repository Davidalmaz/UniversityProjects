CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 1 100 9
32 88 1248 655
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
16 C:\CM60S\BOM.DAT
0 7
32 88 1248 655
143654930 0
0
6 Title:
5 Name:
0
0
0
8
13 Logic Switch~
5 123 244 0 10 11
0 11 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
1 D
-3 -26 4 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
8953 0 0
0
0
13 Logic Switch~
5 121 202 0 1 11
0 12
0
0 0 21360 0
2 0V
-6 -16 8 -8
1 C
-3 -26 4 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
4441 0 0
0
0
13 Logic Switch~
5 125 166 0 1 11
0 13
0
0 0 21360 0
2 0V
-6 -16 8 -8
1 B
-3 -26 4 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
3618 0 0
0
0
13 Logic Switch~
5 124 121 0 10 11
0 14 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
1 A
-3 -26 4 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
6153 0 0
0
0
2 +V
167 539 34 0 1 3
0 9
0
0 0 54256 0
2 5V
-7 -22 7 -14
2 V5
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 0 0
1 V
5394 0 0
0
0
6 74LS47
187 280 184 0 14 29
0 14 13 12 11 15 16 2 3 4
5 6 7 8 17
0
0 0 13040 0
6 74LS47
-21 -60 21 -52
2 U1
-7 -61 7 -53
0
15 DVCC=16;DGND=8;
119 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %14i]
+ [%16bo %1o %2o %3o %4o %5o %6o %14o %7o %8o %9o %10o %11o %12o %13o] %M
0
12 type:digital
5 DIP16
29

0 6 2 1 7 3 5 14 15 9
10 11 12 13 4 6 2 1 7 3
5 14 15 9 10 11 12 13 4 0
65 0 0 512 1 0 0 0
1 U
7734 0 0
0
0
9 CA 7-Seg~
184 447 96 0 18 19
10 8 7 6 5 4 3 2 18 10
0 0 0 2 2 0 0 2 1
0
0 0 21088 0
5 REDCA
16 -41 51 -33
5 DISP1
30 -4 65 4
0
0
32 %D %1 %2 %3 %4 %5 %6 %7 %8 %9 %S
0
0
0
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
88 0 0 512 0 0 0 0
4 DISP
9914 0 0
0
0
9 Resistor~
219 495 46 0 4 5
0 10 9 0 1
0
0 0 880 0
6 0.047k
-20 -14 22 -6
2 R1
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 0 0 0 0
1 R
3747 0 0
0
0
13
7 7 2 0 0 8320 0 7 6 0 0 3
462 132
462 148
318 148
6 8 3 0 0 8320 0 7 6 0 0 3
456 132
456 157
318 157
5 9 4 0 0 8320 0 7 6 0 0 3
450 132
450 166
318 166
4 10 5 0 0 8320 0 7 6 0 0 3
444 132
444 175
318 175
3 11 6 0 0 8320 0 7 6 0 0 3
438 132
438 184
318 184
2 12 7 0 0 8320 0 7 6 0 0 3
432 132
432 193
318 193
1 13 8 0 0 8320 0 7 6 0 0 3
426 132
426 202
318 202
2 1 9 0 0 4224 0 8 5 0 0 3
513 46
539 46
539 43
9 1 10 0 0 8320 0 7 8 0 0 4
447 60
447 50
477 50
477 46
1 4 11 0 0 4224 0 1 6 0 0 6
135 244
239 244
239 173
251 173
251 175
248 175
1 3 12 0 0 8320 0 2 6 0 0 7
133 202
133 205
221 205
221 164
251 164
251 166
248 166
1 2 13 0 0 8320 0 3 6 0 0 5
137 166
137 155
251 155
251 157
248 157
1 1 14 0 0 4240 0 4 6 0 0 6
136 121
236 121
236 146
251 146
251 148
248 148
0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
