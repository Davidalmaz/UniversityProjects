CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 2 100 9
-6 73 757 805
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
16 C:\CM60S\BOM.DAT
0 7
18 585 691 726
160432146 0
0
6 Title:
5 Name:
0
0
0
21
13 Logic Switch~
5 45 43 0 10 11
0 14 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
1 A
-3 -26 4 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
8953 0 0
0
0
13 Logic Switch~
5 43 90 0 10 11
0 13 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
1 B
-3 -26 4 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
4441 0 0
0
0
13 Logic Switch~
5 44 134 0 10 11
0 12 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
1 C
-3 -26 4 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3618 0 0
0
0
13 Logic Switch~
5 44 181 0 10 11
0 11 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
1 D
-3 -26 4 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
6153 0 0
0
0
5 SCOPE
12 550 364 0 1 11
0 3
0
0 0 57584 180
3 SAL
-11 -4 10 4
2 U2
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
0
5394 0 0
0
0
5 SCOPE
12 109 297 0 1 11
0 4
0
0 0 57584 0
4 ENT2
-14 -4 14 4
2 U2
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
0
7734 0 0
0
0
5 SCOPE
12 111 455 0 1 11
0 5
0
0 0 57584 180
4 ENT1
-14 -4 14 4
2 U2
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
0
9914 0 0
0
0
7 Pulser~
4 49 384 0 10 12
0 18 19 4 5 0 0 5 5 3
8
0
0 0 4656 0
0
5 RELOJ
-17 -28 18 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
1 V
3747 0 0
0
0
6 74LS93
109 203 366 0 8 17
0 2 2 4 5 8 7 6 5
0
0 0 13040 0
6 74LS93
-21 -35 21 -27
4 CONT
-14 -36 14 -28
0
15 DVCC=5;DGND=10;
76 %D [%5bi %10bi %1i %2i %3i %4i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o] %M
0
12 type:digital
5 DIP14
17

0 2 3 14 1 11 8 9 12 2
3 14 1 11 8 9 12 0
65 0 0 0 1 0 0 0
1 U
3549 0 0
0
0
10 2-In NAND~
219 402 332 0 3 22
0 8 7 10
0
0 0 112 0
6 74LS00
-14 -24 28 -16
2 A4
0 -34 14 -26
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 2 0
1 U
7931 0 0
0
0
10 2-In NAND~
219 482 335 0 3 22
0 10 9 3
0
0 0 112 0
6 74LS00
-14 -24 28 -16
2 A2
0 -34 14 -26
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 2 0
1 U
9325 0 0
0
0
10 2-In NAND~
219 398 399 0 3 22
0 6 5 9
0
0 0 112 0
6 74LS00
-14 -24 28 -16
2 A3
0 -34 14 -26
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 2 0
1 U
8903 0 0
0
0
10 2-In NAND~
219 490 394 0 3 22
0 20 21 22
0
0 0 112 0
6 74LS00
-14 -24 28 -16
2 A1
0 -34 14 -26
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 512 4 1 2 0
1 U
3834 0 0
0
0
7 Ground~
168 619 340 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3363 0 0
0
0
7 Ground~
168 384 85 0 1 3
0 2
0
0 0 53360 0
0
4 GND2
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
7668 0 0
0
0
10 2-In NAND~
219 251 131 0 3 22
0 23 24 25
0
0 0 112 0
6 74LS00
-14 -24 28 -16
3 A3A
-3 -34 18 -26
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 512 4 1 3 0
1 U
4718 0 0
0
0
10 2-In NAND~
219 163 144 0 3 22
0 12 11 16
0
0 0 112 0
6 74LS00
-14 -24 28 -16
2 A2
0 -34 14 -26
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 3 0
1 U
3874 0 0
0
0
10 2-In NAND~
219 247 80 0 3 22
0 17 16 15
0
0 0 112 0
6 74LS00
-14 -24 28 -16
3 A3C
-3 -34 18 -26
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 3 0
1 U
6671 0 0
0
0
10 2-In NAND~
219 167 77 0 3 22
0 14 13 17
0
0 0 112 0
6 74LS00
-14 -24 28 -16
2 A1
0 -34 14 -26
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 3 0
1 U
3789 0 0
0
0
5 Lamp~
206 607 321 0 2 3
11 3 2
0
0 0 608 0
3 100
-10 -24 11 -16
4 LAMP
-14 -22 14 -14
0
0
11 %D %1 %2 %V
0
0
0
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 L
4871 0 0
0
0
5 Lamp~
206 372 66 0 2 3
11 15 2
0
0 0 608 0
3 100
-10 -24 11 -16
4 LAMP
-14 -22 14 -14
0
0
11 %D %1 %2 %V
0
0
0
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 L
3750 0 0
0
0
24
1 0 3 0 0 4112 0 5 0 0 13 2
548 358
548 334
1 0 4 0 0 4112 0 6 0 0 6 2
109 309
109 375
1 0 5 0 0 4112 0 7 0 0 5 2
109 449
109 384
0 0 5 0 0 8208 0 0 0 5 9 4
153 384
153 403
243 403
243 408
4 4 5 0 0 16 0 8 9 0 0 2
79 384
165 384
3 3 4 0 0 4240 0 9 8 0 0 2
165 375
73 375
2 0 2 0 0 4112 0 9 0 0 8 4
171 366
162 366
162 357
161 357
1 2 2 0 0 12432 0 9 20 0 0 6
171 357
161 357
161 256
633 256
633 334
619 334
2 8 5 0 0 4240 0 12 9 0 0 4
374 408
243 408
243 384
235 384
1 7 6 0 0 8336 0 12 9 0 0 3
374 390
374 375
235 375
2 6 7 0 0 8336 0 10 9 0 0 3
378 341
378 366
235 366
1 5 8 0 0 4240 0 10 9 0 0 4
378 323
243 323
243 357
235 357
3 1 3 0 0 8336 0 11 20 0 0 3
509 335
509 334
595 334
3 2 9 0 0 8336 0 12 11 0 0 4
425 399
448 399
448 344
458 344
3 1 10 0 0 4240 0 10 11 0 0 4
429 332
450 332
450 326
458 326
1 2 2 0 0 16 0 14 20 0 0 2
619 334
619 334
1 2 11 0 0 4224 0 4 17 0 0 4
56 181
131 181
131 153
139 153
1 1 12 0 0 8320 0 3 17 0 0 3
56 134
56 135
139 135
1 2 13 0 0 8320 0 2 19 0 0 3
55 90
55 86
143 86
1 1 14 0 0 4224 0 1 19 0 0 4
57 43
135 43
135 68
143 68
3 1 15 0 0 8320 0 18 21 0 0 3
274 80
274 79
360 79
3 2 16 0 0 8320 0 17 18 0 0 4
190 144
213 144
213 89
223 89
3 1 17 0 0 4224 0 19 18 0 0 4
194 77
215 77
215 71
223 71
1 2 2 0 0 0 0 15 21 0 0 2
384 79
384 79
6
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
377 362 409 386
387 370 411 386
3 CD'
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
381 295 413 319
391 303 415 319
3 AB'
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
445 296 493 320
455 304 495 320
5 AB+CD
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
139 106 171 130
149 114 173 130
3 CD'
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
143 38 175 62
153 46 177 62
3 AB'
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
210 41 258 65
220 49 260 65
5 AB+CD
0
2049 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
788264 1079360 100 100 0 0
0 0 0 0
1 66 162 136
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
12385 0
4 2 2
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
