CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 1 100 9
1 79 585 671
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
16 C:\CM60S\BOM.DAT
0 7
1 79 585 671
143654930 0
0
6 Title:
5 Name:
0
0
0
14
9 2-In AND~
219 344 397 0 3 22
0 4 5 7
0
0 0 624 0
6 74LS08
-21 -24 21 -16
2 BD
-10 -24 4 -16
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 2 0
1 U
8953 0 0
0
0
7 Pulser~
4 55 322 0 10 12
0 12 13 11 14 0 0 5 5 2
7
0
0 0 4656 0
0
3 CLK
-10 -28 11 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
1 V
4441 0 0
0
0
2 +V
167 361 192 0 1 3
0 8
0
0 0 54256 0
2 5V
-7 -22 7 -14
2 V2
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
3618 0 0
0
0
2 +V
167 185 192 0 1 3
0 10
0
0 0 54256 0
2 5V
-7 -22 7 -14
2 V1
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
6153 0 0
0
0
6 74LS76
104 403 268 0 14 29
0 8 8 5 8 8 7 8 6 8
8 4 15 3 9
0
0 0 13040 0
6 74LS76
-21 -60 21 -52
2 U5
-7 -61 7 -53
0
15 DVCC=16;DGND=8;
131 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 4 16 1 2 3 9 12 6 7
8 15 14 11 10 4 16 1 2 3
9 12 6 7 8 15 14 11 10 0
65 0 0 512 1 0 0 0
1 U
5394 0 0
0
0
6 74LS76
104 229 268 0 14 29
0 10 10 11 10 10 9 10 6 10
10 6 16 5 17
0
0 0 13040 0
6 74LS76
-21 -60 21 -52
2 U4
-7 -61 7 -53
0
15 DVCC=16;DGND=8;
131 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 4 16 1 2 3 9 12 6 7
8 15 14 11 10 4 16 1 2 3
9 12 6 7 8 15 14 11 10 0
65 0 0 512 1 0 0 0
1 U
7734 0 0
0
0
7 Ground~
168 294 67 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
9914 0 0
0
0
7 Ground~
168 351 68 0 1 3
0 2
0
0 0 53360 0
0
4 GND2
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3747 0 0
0
0
7 Ground~
168 411 65 0 1 3
0 2
0
0 0 53360 0
0
4 GND3
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3549 0 0
0
0
7 Ground~
168 461 65 0 1 3
0 2
0
0 0 53360 0
0
4 GND4
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
7931 0 0
0
0
5 Lamp~
206 283 48 0 2 3
11 3 2
0
0 0 624 0
3 100
-10 -24 11 -16
1 D
-4 -22 3 -14
0
0
11 %D %1 %2 %V
0
0
0
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 L
9325 0 0
0
0
5 Lamp~
206 339 48 0 2 3
11 4 2
0
0 0 624 0
3 100
-10 -24 11 -16
1 C
-4 -22 3 -14
0
0
11 %D %1 %2 %V
0
0
0
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 L
8903 0 0
0
0
5 Lamp~
206 398 46 0 2 3
11 5 2
0
0 0 624 0
3 100
-10 -24 11 -16
1 B
-4 -22 3 -14
0
0
11 %D %1 %2 %V
0
0
0
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 L
3834 0 0
0
0
5 Lamp~
206 451 46 0 2 3
11 6 2
0
0 0 624 0
3 100
-10 -24 11 -16
1 A
-4 -22 3 -14
0
0
11 %D %1 %2 %V
0
0
0
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 L
3363 0 0
0
0
30
13 1 3 0 0 8320 0 5 11 0 0 5
435 277
448 277
448 97
271 97
271 61
0 1 4 0 0 8192 0 0 12 6 0 5
461 232
461 113
319 113
319 61
327 61
0 1 5 0 0 4224 0 0 13 8 0 5
290 277
290 130
378 130
378 59
386 59
0 1 6 0 0 8320 0 0 14 19 0 5
278 232
278 148
431 148
431 59
439 59
3 6 7 0 0 8320 0 1 5 0 0 6
365 397
369 397
369 327
352 327
352 277
371 277
11 1 4 0 0 12416 0 5 1 0 0 6
435 232
463 232
463 368
312 368
312 388
320 388
0 2 5 0 0 0 0 0 1 8 0 3
302 277
302 406
320 406
13 3 5 0 0 0 0 6 5 0 0 4
261 277
302 277
302 250
365 250
5 0 8 0 0 8192 0 5 0 0 15 3
365 268
365 267
360 267
6 14 9 0 0 12416 0 6 5 0 0 6
197 277
155 277
155 356
449 356
449 286
441 286
4 0 8 0 0 0 0 5 0 0 20 2
365 259
361 259
4 0 10 0 0 4096 0 6 0 0 23 2
191 259
185 259
5 0 10 0 0 0 0 6 0 0 23 2
191 268
185 268
9 0 8 0 0 4096 0 5 0 0 15 2
365 304
335 304
10 0 8 0 0 8320 0 5 0 0 20 4
365 313
335 313
335 267
361 267
9 0 10 0 0 4224 0 6 0 0 17 2
191 304
144 304
0 10 10 0 0 0 0 0 6 23 0 4
185 267
144 267
144 313
191 313
8 0 6 0 0 16 0 5 0 0 19 2
365 295
278 295
11 8 6 0 0 0 0 6 6 0 0 6
261 232
278 232
278 337
183 337
183 295
191 295
7 0 8 0 0 0 0 5 0 0 21 3
371 286
361 286
361 241
2 0 8 0 0 0 0 5 0 0 22 3
371 241
361 241
361 232
1 1 8 0 0 0 0 5 3 0 0 3
371 232
361 232
361 201
7 0 10 0 0 0 0 6 0 0 24 3
197 286
185 286
185 241
2 0 10 0 0 0 0 6 0 0 25 3
197 241
185 241
185 230
1 1 10 0 0 0 0 4 6 0 0 3
185 201
185 232
197 232
1 2 2 0 0 4224 0 10 14 0 0 2
461 59
463 59
1 2 2 0 0 0 0 9 13 0 0 2
411 59
410 59
1 2 2 0 0 0 0 8 12 0 0 2
351 62
351 61
1 2 2 0 0 0 0 7 11 0 0 2
294 61
295 61
3 3 11 0 0 24704 0 2 6 0 0 7
79 313
79 316
78 316
78 314
109 314
109 250
191 250
0
0
2049 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
1967336 1079360 100 100 0 0
0 0 0 0
2 74 163 144
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
12385 0
4 0.05 2
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
