CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
240 0 30 100 9
871 90 1575 807
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
16 C:\CM60S\BOM.DAT
0 7
871 90 1575 807
143654930 0
0
6 Title:
5 Name:
0
0
0
29
13 Logic Switch~
5 341 894 0 1 11
0 4
0
0 0 21360 0
2 0V
-6 -16 8 -8
1 B
-3 -26 4 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
8953 0 0
0
0
13 Logic Switch~
5 342 825 0 10 11
0 5 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -18 8 -10
1 A
-2 -30 5 -22
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
4441 0 0
0
0
13 Logic Switch~
5 341 670 0 10 11
0 8 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -18 8 -10
1 A
-2 -30 5 -22
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
3618 0 0
0
0
13 Logic Switch~
5 340 739 0 1 11
0 7
0
0 0 21360 0
2 0V
-6 -16 8 -8
1 B
-3 -26 4 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
6153 0 0
0
0
13 Logic Switch~
5 336 594 0 1 11
0 10
0
0 0 21360 0
2 0V
-6 -16 8 -8
1 B
-3 -26 4 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5394 0 0
0
0
13 Logic Switch~
5 337 525 0 10 11
0 11 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -18 8 -10
1 A
-2 -30 5 -22
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
7734 0 0
0
0
13 Logic Switch~
5 332 422 0 1 11
0 13
0
0 0 21360 0
2 0V
-6 -16 8 -8
1 A
-3 -26 4 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
9914 0 0
0
0
13 Logic Switch~
5 328 253 0 10 11
0 16 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -18 8 -10
1 A
-2 -30 5 -22
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
3747 0 0
0
0
13 Logic Switch~
5 327 322 0 10 11
0 15 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
1 B
-3 -26 4 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
3549 0 0
0
0
13 Logic Switch~
5 323 156 0 10 11
0 18 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
1 B
-3 -26 4 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
7931 0 0
0
0
13 Logic Switch~
5 324 87 0 10 11
0 19 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -18 8 -10
1 A
-2 -30 5 -22
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
9325 0 0
0
0
7 Ground~
168 731 866 0 1 3
0 2
0
0 0 53360 0
0
4 GND5
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
8903 0 0
0
0
9 2-In XOR~
219 503 857 0 3 22
0 5 4 3
0
0 0 624 0
6 74LS86
-21 -24 21 -16
3 XOR
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 4 0
1 U
3834 0 0
0
0
7 Ground~
168 727 709 0 1 3
0 2
0
0 0 53360 0
0
4 GND3
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3363 0 0
0
0
8 2-In OR~
219 499 701 0 3 22
0 8 7 6
0
0 0 624 0
6 74LS32
-21 -24 21 -16
2 OR
0 -25 14 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0
65 0 0 0 4 1 3 0
1 U
7668 0 0
0
0
7 Ground~
168 728 564 0 1 3
0 2
0
0 0 53360 0
0
4 GND6
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
4718 0 0
0
0
9 2-In AND~
219 500 555 0 3 22
0 11 10 9
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 AND
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 5 0
1 U
3874 0 0
0
0
7 Ground~
168 725 431 0 1 3
0 2
0
0 0 53360 0
0
4 GND2
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
6671 0 0
0
0
9 Inverter~
13 496 422 0 2 22
0 13 12
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 NOT
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
15

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0
65 0 0 0 6 1 2 0
1 U
3789 0 0
0
0
7 Ground~
168 722 289 0 1 3
0 2
0
0 0 53360 0
0
4 GND7
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
4871 0 0
0
0
9 2-In NOR~
219 485 283 0 3 22
0 16 15 14
0
0 0 112 0
6 74LS02
-21 -24 21 -16
1 N
-4 -34 3 -26
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0
65 0 0 0 4 2 6 0
1 U
3750 0 0
0
0
7 Ground~
168 716 124 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
8778 0 0
0
0
10 2-In NAND~
219 492 118 0 3 22
0 19 18 17
0
0 0 624 0
6 74LS00
-14 -24 28 -16
4 NAND
-16 -30 12 -22
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 1138729552
65 0 0 0 4 1 1 0
1 U
538 0 0
0
0
5 Lamp~
206 719 845 0 2 3
11 3 2
0
0 0 608 0
3 100
-10 -24 11 -16
2 S6
-7 -22 7 -14
0
0
11 %D %1 %2 %V
0
0
0
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 L
6843 0 0
0
0
5 Lamp~
206 715 688 0 2 3
11 6 2
0
0 0 608 0
3 100
-10 -24 11 -16
2 S5
-7 -22 7 -14
0
0
11 %D %1 %2 %V
0
0
0
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 L
3136 0 0
0
0
5 Lamp~
206 716 543 0 2 3
11 9 2
0
0 0 608 0
3 100
-10 -24 11 -16
2 S4
-7 -22 7 -14
0
0
11 %D %1 %2 %V
0
0
0
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 L
5950 0 0
0
0
5 Lamp~
206 713 410 0 2 3
11 12 2
0
0 0 608 0
3 100
-10 -24 11 -16
2 S3
-7 -22 7 -14
0
0
11 %D %1 %2 %V
0
0
0
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 L
5670 0 0
0
0
5 Lamp~
206 710 268 0 2 3
11 14 2
0
0 0 608 0
3 100
-10 -24 11 -16
2 S2
-7 -22 7 -14
0
0
11 %D %1 %2 %V
0
0
0
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 L
6828 0 0
0
0
5 Lamp~
206 704 103 0 2 3
11 17 2
0
0 0 608 0
3 100
-10 -24 11 -16
2 S1
-7 -22 7 -14
0
0
11 %D %1 %2 %V
0
0
0
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 L
6735 0 0
0
0
23
1 2 2 0 0 4224 0 12 24 0 0 4
731 860
731 856
731 856
731 858
3 1 3 0 0 8320 0 13 24 0 0 4
536 857
536 857
707 857
707 858
1 2 4 0 0 4224 0 1 13 0 0 3
353 894
487 894
487 866
1 1 5 0 0 8320 0 2 13 0 0 4
354 825
354 828
487 828
487 848
1 2 2 0 0 0 0 14 25 0 0 4
727 703
727 699
727 699
727 701
3 1 6 0 0 8320 0 15 25 0 0 4
532 701
532 700
703 700
703 701
1 2 7 0 0 4224 0 4 15 0 0 3
352 739
486 739
486 710
1 1 8 0 0 8320 0 3 15 0 0 4
353 670
353 673
486 673
486 692
1 2 2 0 0 0 0 16 26 0 0 4
728 558
728 554
728 554
728 556
3 1 9 0 0 4224 0 17 26 0 0 3
521 555
704 555
704 556
1 2 10 0 0 4224 0 5 17 0 0 3
348 594
476 594
476 564
1 1 11 0 0 4224 0 6 17 0 0 3
349 525
476 525
476 546
1 2 2 0 0 0 0 18 27 0 0 4
725 425
725 421
725 421
725 423
2 1 12 0 0 4224 0 19 27 0 0 3
517 422
701 422
701 423
1 1 13 0 0 4224 0 7 19 0 0 2
344 422
481 422
1 2 2 0 0 0 0 20 28 0 0 2
722 283
722 281
3 1 14 0 0 4224 0 21 28 0 0 4
524 283
700 283
700 281
698 281
1 2 15 0 0 4224 0 9 21 0 0 3
339 322
472 322
472 292
1 1 16 0 0 4224 0 8 21 0 0 3
340 253
472 253
472 274
1 2 2 0 0 0 0 22 29 0 0 2
716 118
716 116
3 1 17 0 0 4224 0 23 29 0 0 4
519 118
694 118
694 116
692 116
1 2 18 0 0 4224 0 10 23 0 0 3
335 156
468 156
468 127
1 1 19 0 0 4224 0 11 23 0 0 3
336 87
468 87
468 109
11
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
468 242 500 266
478 250 502 266
3 NOR
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 4
240 695 280 719
248 703 280 719
4 7432
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 4
234 402 274 426
244 410 276 426
4 7404
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 4
245 844 285 868
255 852 287 868
4 7486
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 4
239 542 279 566
249 550 281 566
4 7408
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 4
229 278 269 302
239 286 271 302
4 7402
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 4
224 103 264 127
234 111 266 127
4 7400
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 8
283 12 355 36
293 20 357 36
8 ENTRADAS
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 18
425 14 577 38
435 21 579 37
18 COMPUERTAS L�GICAS
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 6
670 15 726 39
680 23 728 39
6 SALIDA
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
233 14 257 38
241 22 257 38
2 CI
0
2049 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
