CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 90 30 100 9
32 88 1248 655
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
16 C:\CM60S\BOM.DAT
0 7
32 88 1248 655
143654930 0
0
6 Title:
5 Name:
0
0
0
15
13 Logic Switch~
5 253 294 0 1 11
0 11
0
0 0 21360 0
2 0V
-6 -16 8 -8
1 D
-3 -26 4 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
8953 0 0
0
0
13 Logic Switch~
5 254 213 0 1 11
0 9
0
0 0 21360 0
2 0V
-6 -16 8 -8
1 C
-3 -26 4 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
4441 0 0
0
0
13 Logic Switch~
5 253 133 0 1 11
0 7
0
0 0 21360 0
2 0V
-6 -16 8 -8
1 B
-3 -26 4 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3618 0 0
0
0
10 2-In NAND~
219 414 507 0 3 22
0 7 3 4
0
0 0 624 0
6 74LS00
-14 -24 28 -16
3 U3B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 3 0
1 U
6153 0 0
0
0
10 2-In NAND~
219 409 459 0 3 22
0 6 3 5
0
0 0 624 0
6 74LS00
-14 -24 28 -16
3 U3A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 3 0
1 U
5394 0 0
0
0
10 2-In NAND~
219 522 455 0 3 22
0 5 4 8
0
0 0 624 0
6 74LS00
-14 -24 28 -16
3 U2D
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 2 0
1 U
7734 0 0
0
0
7 Ground~
168 596 470 0 1 3
0 2
0
0 0 53360 0
0
4 GND2
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
9914 0 0
0
0
10 2-In NAND~
219 336 450 0 3 22
0 9 9 6
0
0 0 624 0
6 74LS00
-14 -24 28 -16
3 U2B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 2 0
1 U
3747 0 0
0
0
10 2-In NAND~
219 505 209 0 3 22
0 10 3 13
0
0 0 624 0
6 74LS00
-14 -24 28 -16
3 U1D
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 1 0
1 U
3549 0 0
0
0
10 2-In NAND~
219 337 284 0 3 22
0 11 11 3
0
0 0 624 0
6 74LS00
-14 -24 28 -16
3 U1C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 1 0
1 U
7931 0 0
0
0
10 2-In NAND~
219 396 171 0 3 22
0 12 9 10
0
0 0 624 0
6 74LS00
-14 -24 28 -16
3 U1B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 1 0
1 U
9325 0 0
0
0
10 2-In NAND~
219 332 127 0 3 22
0 7 7 12
0
0 0 624 0
6 74LS00
-14 -24 28 -16
3 U1A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 1 0
1 U
8903 0 0
0
0
7 Ground~
168 582 219 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3834 0 0
0
0
5 Lamp~
206 585 443 0 2 3
11 8 2
0
0 0 624 0
3 100
-10 -24 11 -16
2 L2
-7 -22 7 -14
0
0
11 %D %1 %2 %V
0
0
0
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 L
3363 0 0
0
0
5 Lamp~
206 569 195 0 2 3
11 13 2
0
0 0 624 0
3 100
-10 -24 11 -16
2 L1
-7 -22 7 -14
0
0
11 %D %1 %2 %V
0
0
0
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 L
7668 0 0
0
0
20
3 2 3 0 0 8336 0 10 4 0 0 4
364 284
368 284
368 516
390 516
3 2 4 0 0 4224 0 4 6 0 0 3
441 507
498 507
498 464
3 1 5 0 0 8320 0 5 6 0 0 3
436 459
436 446
498 446
3 1 6 0 0 4224 0 8 5 0 0 2
363 450
385 450
0 2 3 0 0 128 0 0 5 1 0 3
376 516
376 468
385 468
0 1 7 0 0 4224 0 0 4 18 0 3
281 133
281 498
390 498
3 1 8 0 0 8320 0 6 14 0 0 3
549 455
549 456
573 456
0 2 9 0 0 8192 0 0 8 9 0 3
291 446
291 459
312 459
0 1 9 0 0 4224 0 0 8 16 0 5
291 213
291 446
291 446
291 441
312 441
1 2 2 0 0 4224 0 7 14 0 0 3
596 464
596 456
597 456
3 1 10 0 0 4224 0 11 9 0 0 4
423 171
473 171
473 200
481 200
3 2 3 0 0 128 0 10 9 0 0 4
364 284
473 284
473 218
481 218
0 1 11 0 0 4096 0 0 10 14 0 3
302 294
302 275
313 275
1 2 11 0 0 4224 0 1 10 0 0 4
265 294
305 294
305 293
313 293
3 1 12 0 0 8320 0 12 11 0 0 4
359 127
364 127
364 162
372 162
1 2 9 0 0 0 0 2 11 0 0 4
266 213
364 213
364 180
372 180
0 2 7 0 0 0 0 0 12 18 0 3
299 133
299 136
308 136
1 1 7 0 0 0 0 3 12 0 0 4
265 133
300 133
300 118
308 118
3 1 13 0 0 12416 0 9 15 0 0 4
532 209
533 209
533 208
557 208
1 2 2 0 0 0 0 13 15 0 0 3
582 213
582 208
581 208
0
0
2049 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
592174 1079360 100 100 0 0
0 0 0 0
1 66 162 136
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
12385 0
4 0.5 2
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
