CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 5 100 9
0 71 1536 824
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
16 C:\CM60S\BOM.DAT
0 7
0 71 1536 824
143654930 0
0
6 Title:
5 Name:
0
0
0
7
13 Logic Switch~
5 113 141 0 1 11
0 3
0
0 0 21344 0
2 0V
-7 -15 7 -7
2 V2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
8953 0 0
0
0
10 2-In NAND~
219 236 131 0 3 22
0 5 6 7
0
0 0 608 0
6 74LS00
-14 -24 28 -16
4 NAND
-7 -34 21 -26
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 512 4 4 1 0
1 U
4441 0 0
0
0
10 2-In NAND~
219 381 134 0 3 22
0 8 3 4
0
0 0 608 0
6 74LS00
-14 -24 28 -16
4 NAND
-7 -34 21 -26
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 512 4 3 1 0
1 U
3618 0 0
0
0
10 2-In NAND~
219 236 261 0 3 22
0 9 10 11
0
0 0 608 0
6 74LS00
-14 -24 28 -16
4 NAND
-7 -34 21 -26
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 512 4 2 1 0
1 U
6153 0 0
0
0
10 2-In NAND~
219 385 267 0 3 22
0 12 13 14
0
0 0 608 0
6 74LS00
-14 -24 28 -16
4 NAND
-7 -34 21 -26
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 512 4 1 1 0
1 U
5394 0 0
0
0
7 Ground~
168 816 141 0 1 3
0 2
0
0 0 53344 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
7734 0 0
0
0
5 Lamp~
206 589 121 0 2 3
11 4 2
0
0 0 624 0
3 100
-10 -24 11 -16
4 LAMP
-14 -22 14 -14
0
0
11 %D %1 %2 %V
0
0
0
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 L
9914 0 0
0
0
3
1 2 3 0 0 4224 0 1 3 0 0 6
125 141
208 141
208 151
288 151
288 143
357 143
3 1 4 0 0 4224 0 3 7 0 0 2
408 134
577 134
1 2 2 0 0 4224 0 6 7 0 0 3
816 135
601 135
601 134
0
0
2049 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
1117004 1079360 100 100 0 0
0 0 0 0
1 66 162 136
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
12385 0
4 0.5 2
1
383 131
0 4 0 0 1	0 2 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
