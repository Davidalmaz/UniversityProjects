CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 910 30 100 9
3 80 659 824
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
18 C:\CM50_32\BOM.DAT
0 7
3 80 659 824
143654930 0
0
6 Title:
5 Name:
0
0
0
47
13 Logic Switch~
5 132 992 0 1 11
0 8
0
0 0 21360 0
2 0V
-7 -15 7 -7
2 V7
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
8953 0 0
0
0
13 Logic Switch~
5 131 1078 0 1 11
0 7
0
0 0 21360 0
2 0V
-7 -15 7 -7
2 V8
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
4441 0 0
0
0
13 Logic Switch~
5 114 1299 0 10 11
0 9 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-7 -15 7 -7
1 B
-2 -26 5 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3618 0 0
0
0
13 Logic Switch~
5 115 1213 0 10 11
0 10 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-7 -15 7 -7
1 A
-2 -26 5 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
6153 0 0
0
0
13 Logic Switch~
5 103 741 0 10 11
0 19 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-7 -15 7 -7
2 V6
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5394 0 0
0
0
13 Logic Switch~
5 104 810 0 10 11
0 15 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-7 -15 7 -7
2 V5
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
7734 0 0
0
0
13 Logic Switch~
5 107 521 0 1 11
0 23
0
0 0 21360 0
2 0V
-7 -15 7 -7
2 V3
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
9914 0 0
0
0
13 Logic Switch~
5 105 594 0 1 11
0 22
0
0 0 21360 0
2 0V
-7 -15 7 -7
2 V4
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3747 0 0
0
0
13 Logic Switch~
5 94 286 0 1 11
0 29
0
0 0 21360 0
2 0V
-7 -15 7 -7
2 V1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3549 0 0
0
0
13 Logic Switch~
5 93 341 0 1 11
0 28
0
0 0 21360 0
2 0V
-7 -15 7 -7
2 V2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
7931 0 0
0
0
13 Logic Switch~
5 109 108 0 10 11
0 30 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-7 -15 7 -7
2 V1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
9325 0 0
0
0
10 2-In NAND~
219 255 982 0 3 22
0 6 8 5
0
0 0 624 0
6 74LS00
-14 -24 28 -16
5 NAN3A
-10 -34 25 -26
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 5 0
1 U
8903 0 0
0
0
10 2-In NAND~
219 335 985 0 3 22
0 5 4 3
0
0 0 624 0
6 74LS00
-14 -24 28 -16
5 NAN3B
-10 -34 25 -26
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 5 0
1 U
3834 0 0
0
0
10 2-In NAND~
219 251 1049 0 3 22
0 8 7 6
0
0 0 624 0
6 74LS00
-14 -24 28 -16
5 NAN3C
-10 -33 25 -25
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 5 0
1 U
3363 0 0
0
0
10 2-In NAND~
219 329 1049 0 3 22
0 6 7 4
0
0 0 624 0
6 74LS00
-14 -24 28 -16
5 NAN3D
-10 -34 25 -26
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 5 0
1 U
7668 0 0
0
0
7 Ground~
168 472 990 0 1 3
0 2
0
0 0 53360 0
0
4 GND5
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
4718 0 0
0
0
10 2-In NAND~
219 169 1239 0 3 22
0 10 9 11
0
0 0 624 0
6 74LS00
-14 -24 28 -16
5 NAN4A
-10 -33 25 -25
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 6 0
1 U
3874 0 0
0
0
10 2-In NAND~
219 219 1322 0 3 22
0 11 9 12
0
0 0 624 0
6 74LS00
-14 -24 28 -16
5 NAN4B
-10 -34 25 -26
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 6 0
1 U
6671 0 0
0
0
10 2-In NAND~
219 433 1255 0 3 22
0 13 12 14
0
0 0 624 0
6 74LS00
-14 -24 28 -16
5 NAN4C
-10 -34 25 -26
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 6 0
1 U
3789 0 0
0
0
10 2-In NAND~
219 226 1169 0 3 22
0 10 11 13
0
0 0 624 0
6 74LS00
-14 -24 28 -16
5 NAN4D
-10 -34 25 -26
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 6 0
1 U
4871 0 0
0
0
7 Ground~
168 523 1261 0 1 3
0 2
0
0 0 53360 0
0
4 GND6
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3750 0 0
0
0
10 2-In NAND~
219 208 732 0 3 22
0 32 19 20
0
0 0 624 0
6 74LS00
-14 -24 28 -16
5 NAN2D
-10 -34 25 -26
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 512 4 4 4 0
1 U
8778 0 0
0
0
10 2-In NAND~
219 396 737 0 3 22
0 20 18 17
0
0 0 624 0
6 74LS00
-14 -24 28 -16
5 NAN2C
-10 -34 25 -26
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 4 0
1 U
538 0 0
0
0
10 2-In NAND~
219 209 803 0 3 22
0 33 15 18
0
0 0 624 0
6 74LS00
-14 -24 28 -16
5 NAN2B
-10 -34 25 -26
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 512 4 2 4 0
1 U
6843 0 0
0
0
10 2-In NAND~
219 448 818 0 3 22
0 17 34 16
0
0 0 624 0
6 74LS00
-14 -24 28 -16
5 NAN2A
-10 -34 25 -26
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 512 4 1 4 0
1 U
3136 0 0
0
0
7 Ground~
168 602 831 0 1 3
0 2
0
0 0 53360 0
0
4 GND4
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
5950 0 0
0
0
10 2-In NAND~
219 230 511 0 3 22
0 35 23 24
0
0 0 624 0
6 74LS00
-14 -24 28 -16
5 NAN1D
-10 -34 25 -26
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 512 4 4 3 0
1 U
5670 0 0
0
0
10 2-In NAND~
219 478 514 0 3 22
0 24 21 25
0
0 0 624 0
6 74LS00
-14 -24 28 -16
5 NAN1C
-10 -34 25 -26
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 3 0
1 U
6828 0 0
0
0
10 2-In NAND~
219 236 585 0 3 22
0 36 22 21
0
0 0 624 0
6 74LS00
-14 -24 28 -16
5 NAN1B
-10 -34 25 -26
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 512 4 2 3 0
1 U
6735 0 0
0
0
10 2-In NAND~
219 483 575 0 3 22
0 37 38 39
0
0 0 624 0
6 74LS00
-14 -24 28 -16
5 NAN1A
-10 -35 25 -27
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 512 4 1 3 0
1 U
8365 0 0
0
0
7 Ground~
168 586 520 0 1 3
0 2
0
0 0 53360 0
0
4 GND3
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
4132 0 0
0
0
7 Ground~
168 598 316 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
4551 0 0
0
0
10 2-In NAND~
219 353 381 0 3 22
0 40 41 42
0
0 0 624 0
6 74LS00
-14 -24 28 -16
4 NAND
-7 -34 21 -26
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 512 4 4 2 0
1 U
3635 0 0
0
0
10 2-In NAND~
219 220 377 0 3 22
0 43 44 45
0
0 0 624 0
6 74LS00
-14 -24 28 -16
4 NAND
-7 -34 21 -26
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 512 4 3 2 0
1 U
3973 0 0
0
0
10 2-In NAND~
219 389 305 0 3 22
0 26 46 27
0
0 0 624 0
6 74LS00
-14 -24 28 -16
4 NAND
-7 -34 21 -26
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 512 4 2 2 0
1 U
3851 0 0
0
0
10 2-In NAND~
219 221 306 0 3 22
0 29 28 26
0
0 0 624 0
6 74LS00
-14 -24 28 -16
4 NAND
-6 -33 22 -25
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 2 0
1 U
8383 0 0
0
0
7 Ground~
168 590 108 0 1 3
0 2
0
0 0 53360 0
0
4 GND2
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
9334 0 0
0
0
10 2-In NAND~
219 371 166 0 3 22
0 47 48 49
0
0 0 624 0
6 74LS00
-14 -24 28 -16
4 NAND
-7 -34 21 -26
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 512 4 4 1 0
1 U
7471 0 0
0
0
10 2-In NAND~
219 232 170 0 3 22
0 50 51 52
0
0 0 624 0
6 74LS00
-14 -24 28 -16
4 NANC
-7 -34 21 -26
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 512 4 3 1 0
1 U
3334 0 0
0
0
10 2-In NAND~
219 377 101 0 3 22
0 53 30 31
0
0 0 624 0
6 74LS00
-14 -24 28 -16
4 NANB
-7 -34 21 -26
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 512 4 2 1 0
1 U
3559 0 0
0
0
10 2-In NAND~
219 232 98 0 3 22
0 54 55 56
0
0 0 624 0
6 74LS00
-14 -24 28 -16
4 NANA
-7 -34 21 -26
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 512 4 1 1 0
1 U
984 0 0
0
0
5 Lamp~
206 460 971 0 2 3
11 3 2
0
0 0 608 0
3 100
-10 -24 11 -16
5 LAMP4
-17 -22 18 -14
0
0
11 %D %1 %2 %V
0
0
0
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 L
7557 0 0
0
0
5 Lamp~
206 511 1242 0 2 3
11 14 2
0
0 0 608 0
3 100
-10 -24 11 -16
5 LAMP5
-17 -22 18 -14
0
0
11 %D %1 %2 %V
0
0
0
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 L
3146 0 0
0
0
5 Lamp~
206 541 809 0 2 3
11 16 2
0
0 0 608 0
3 100
-10 -24 11 -16
5 LAMP3
-17 -22 18 -14
0
0
11 %D %1 %2 %V
0
0
0
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 L
5687 0 0
0
0
5 Lamp~
206 540 501 0 2 3
11 25 2
0
0 0 608 0
3 100
-10 -24 11 -16
5 LAMP2
-17 -22 18 -14
0
0
11 %D %1 %2 %V
0
0
0
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 L
7939 0 0
0
0
5 Lamp~
206 489 292 0 2 3
11 27 2
0
0 0 608 0
3 100
-10 -24 11 -16
5 LAMP1
-17 -22 18 -14
0
0
11 %D %1 %2 %V
0
0
0
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 L
3308 0 0
0
0
5 Lamp~
206 478 88 0 2 3
11 31 2
0
0 0 608 0
3 100
-10 -24 11 -16
4 LAMP
-14 -22 14 -14
0
0
11 %D %1 %2 %V
0
0
0
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 L
3408 0 0
0
0
41
3 1 3 0 0 8320 0 13 42 0 0 3
362 985
362 984
448 984
3 2 4 0 0 8320 0 15 13 0 0 6
356 1049
356 1024
313 1024
313 997
311 997
311 994
3 1 5 0 0 4224 0 12 13 0 0 3
282 982
311 982
311 976
0 1 6 0 0 12416 0 0 12 5 0 5
290 1040
290 1096
210 1096
210 973
231 973
3 1 6 0 0 0 0 14 15 0 0 3
278 1049
278 1040
305 1040
0 2 7 0 0 4096 0 0 15 9 0 3
227 1078
305 1078
305 1058
0 2 8 0 0 8192 0 0 12 8 0 3
191 992
191 991
231 991
1 1 8 0 0 8320 0 1 14 0 0 4
144 992
191 992
191 1040
227 1040
1 2 7 0 0 4224 0 2 14 0 0 3
143 1078
227 1078
227 1058
1 2 2 0 0 0 0 16 42 0 0 2
472 984
472 984
1 2 9 0 0 4096 0 3 17 0 0 3
126 1299
126 1248
145 1248
1 1 10 0 0 8192 0 4 17 0 0 3
127 1213
127 1230
145 1230
0 2 11 0 0 4096 0 0 20 14 0 3
194 1241
194 1178
202 1178
3 1 11 0 0 8320 0 17 18 0 0 4
196 1239
194 1239
194 1313
195 1313
1 2 9 0 0 8320 0 3 18 0 0 3
126 1299
126 1331
195 1331
1 1 10 0 0 8320 0 4 20 0 0 3
127 1213
127 1160
202 1160
3 2 12 0 0 4224 0 18 19 0 0 4
246 1322
401 1322
401 1264
409 1264
3 1 13 0 0 4224 0 20 19 0 0 4
253 1169
401 1169
401 1246
409 1246
3 1 14 0 0 4224 0 19 43 0 0 2
460 1255
499 1255
1 2 2 0 0 0 0 21 43 0 0 2
523 1255
523 1255
2 1 2 0 0 4096 0 44 26 0 0 3
553 822
602 822
602 825
1 2 15 0 0 8320 0 6 24 0 0 3
116 810
116 812
185 812
3 1 16 0 0 4224 0 25 44 0 0 3
475 818
529 818
529 822
3 1 17 0 0 4224 0 23 25 0 0 4
423 737
423 808
424 808
424 809
3 2 18 0 0 12416 0 24 23 0 0 4
236 803
264 803
264 746
372 746
1 2 19 0 0 4224 0 5 22 0 0 2
115 741
184 741
3 1 20 0 0 4224 0 22 23 0 0 3
235 732
372 732
372 728
3 2 21 0 0 4224 0 29 28 0 0 4
263 585
446 585
446 523
454 523
1 2 22 0 0 4224 0 8 29 0 0 2
117 594
212 594
1 2 23 0 0 8320 0 7 27 0 0 3
119 521
119 520
206 520
3 1 24 0 0 4224 0 27 28 0 0 3
257 511
454 511
454 505
1 2 2 0 0 0 0 31 45 0 0 2
586 514
552 514
3 1 25 0 0 4224 0 28 45 0 0 2
505 514
528 514
2 1 2 0 0 4096 0 46 32 0 0 3
501 305
598 305
598 310
3 1 26 0 0 4224 0 36 35 0 0 4
248 306
357 306
357 296
365 296
3 1 27 0 0 4224 0 35 46 0 0 2
416 305
477 305
1 2 28 0 0 4224 0 10 36 0 0 4
105 341
189 341
189 315
197 315
1 1 29 0 0 4224 0 9 36 0 0 4
106 286
189 286
189 297
197 297
1 2 30 0 0 4224 0 11 40 0 0 6
121 108
204 108
204 118
284 118
284 110
353 110
3 1 31 0 0 4224 0 40 47 0 0 2
404 101
466 101
1 2 2 0 0 4224 0 37 47 0 0 3
590 102
490 102
490 101
5
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
92 884 124 908
102 892 126 908
3 XOR
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
93 448 117 472
103 456 119 472
2 OR
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
80 209 112 233
90 217 114 233
3 AND
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
91 29 123 53
101 37 125 53
3 NOT
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
86 648 118 672
96 656 120 672
3 NOR
0
2049 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
