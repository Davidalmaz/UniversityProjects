CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 390 30 100 9
32 88 1248 655
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
16 C:\CM60S\BOM.DAT
0 7
32 88 1248 655
143654930 0
0
6 Title:
5 Name:
0
0
0
21
13 Logic Switch~
5 261 539 0 10 11
0 9 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 X1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
8953 0 0
0
0
13 Logic Switch~
5 249 673 0 10 11
0 8 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 Y1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
4441 0 0
0
0
13 Logic Switch~
5 242 762 0 10 11
0 7 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 Z1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
3618 0 0
0
0
13 Logic Switch~
5 202 337 0 1 11
0 14
0
0 0 21360 0
2 0V
-6 -16 8 -8
1 Z
-3 -26 4 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
6153 0 0
0
0
13 Logic Switch~
5 209 248 0 1 11
0 18
0
0 0 21360 0
2 0V
-6 -16 8 -8
1 Y
-3 -26 4 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
5394 0 0
0
0
13 Logic Switch~
5 221 114 0 1 11
0 16
0
0 0 21360 0
2 0V
-6 -16 8 -8
1 X
-3 -26 4 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
7734 0 0
0
0
7 Ground~
168 650 627 0 1 3
0 2
0
0 0 53360 0
0
4 GND2
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
9914 0 0
0
0
10 2-In NAND~
219 601 619 0 3 22
0 5 4 3
0
0 0 624 0
6 74LS00
-14 -24 28 -16
3 U4A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 4 0
1 U
3747 0 0
0
0
10 2-In NAND~
219 485 687 0 3 22
0 8 7 4
0
0 0 624 0
6 74LS00
-14 -24 28 -16
3 U3D
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 3 0
1 U
3549 0 0
0
0
10 2-In NAND~
219 448 551 0 3 22
0 9 6 5
0
0 0 624 0
6 74LS00
-14 -24 28 -16
3 U3C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 3 0
1 U
7931 0 0
0
0
10 2-In NAND~
219 398 668 0 3 22
0 8 8 6
0
0 0 624 0
6 74LS00
-14 -24 28 -16
3 U3B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 3 0
1 U
9325 0 0
0
0
7 Ground~
168 780 241 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
8903 0 0
0
0
10 2-In NAND~
219 512 282 0 3 22
0 16 14 11
0
0 0 624 0
6 74LS00
-14 -24 28 -16
3 U1D
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 1 0
1 U
3834 0 0
0
0
5 4023~
219 732 234 0 4 22
0 13 12 11 10
0
0 0 624 0
4 4023
-14 -28 14 -20
3 U2C
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
17

0 11 12 13 10 3 4 5 6 1
2 8 9 11 12 13 10 0
65 0 0 0 3 3 2 0
1 U
3363 0 0
0
0
5 4023~
219 531 164 0 4 22
0 19 18 14 12
0
0 0 624 0
4 4023
-14 -28 14 -20
3 U2B
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
17

0 1 2 8 9 3 4 5 6 1
2 8 9 11 12 13 10 0
65 0 0 0 3 2 2 0
1 U
7668 0 0
0
0
5 4023~
219 544 93 0 4 22
0 16 17 15 13
0
0 0 624 0
4 4023
-14 -28 14 -20
3 U2A
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
17

0 3 4 5 6 3 4 5 6 1
2 8 9 11 12 13 10 0
65 0 0 0 3 1 2 0
1 U
4718 0 0
0
0
10 2-In NAND~
219 353 328 0 3 22
0 14 14 15
0
0 0 624 0
6 74LS00
-14 -24 28 -16
3 U1C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 1 0
1 U
3874 0 0
0
0
10 2-In NAND~
219 358 243 0 3 22
0 18 18 17
0
0 0 624 0
6 74LS00
-14 -24 28 -16
3 U1B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 1 0
1 U
6671 0 0
0
0
10 2-In NAND~
219 354 136 0 3 22
0 16 16 19
0
0 0 624 0
6 74LS00
-14 -24 28 -16
3 U1A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 1 0
1 U
3789 0 0
0
0
5 Lamp~
206 639 607 0 2 3
11 3 2
0
0 0 608 0
3 100
-10 -24 11 -16
2 L2
-7 -22 7 -14
0
0
11 %D %1 %2 %V
0
0
0
5

0 1 2 1 2 0
82 0 0 0 0 0 0 0
1 L
4871 0 0
0
0
5 Lamp~
206 769 221 0 2 3
11 10 2
0
0 0 608 0
3 100
-10 -24 11 -16
2 L1
-7 -22 7 -14
0
0
11 %D %1 %2 %V
0
0
0
5

0 1 2 1 2 0
82 0 0 0 0 0 0 0
1 L
3750 0 0
0
0
29
1 2 2 0 0 4240 0 7 20 0 0 3
650 621
650 620
651 620
1 3 3 0 0 4240 0 20 8 0 0 3
627 620
628 620
628 619
3 2 4 0 0 8320 0 9 8 0 0 4
512 687
569 687
569 628
577 628
3 1 5 0 0 4224 0 10 8 0 0 4
475 551
569 551
569 610
577 610
3 2 6 0 0 8320 0 11 10 0 0 6
425 668
429 668
429 570
419 570
419 560
424 560
1 2 7 0 0 4224 0 3 9 0 0 4
254 762
453 762
453 696
461 696
0 1 8 0 0 8320 0 0 9 10 0 5
339 673
339 688
453 688
453 678
461 678
1 1 9 0 0 4224 0 1 10 0 0 4
273 539
416 539
416 542
424 542
0 2 8 0 0 0 0 0 11 10 0 3
366 673
366 677
374 677
1 1 8 0 0 0 0 2 11 0 0 4
261 673
366 673
366 659
374 659
1 2 2 0 0 128 0 12 21 0 0 3
780 235
780 234
781 234
1 4 10 0 0 4224 0 21 14 0 0 2
757 234
759 234
3 3 11 0 0 4224 0 13 14 0 0 4
539 282
700 282
700 243
708 243
4 2 12 0 0 8320 0 15 14 0 0 3
558 164
558 234
708 234
4 1 13 0 0 8320 0 16 14 0 0 4
571 93
700 93
700 225
708 225
0 3 14 0 0 4096 0 0 15 20 0 3
450 291
450 173
507 173
3 3 15 0 0 8320 0 17 16 0 0 4
380 328
417 328
417 102
520 102
2 0 14 0 0 0 0 17 0 0 19 4
329 337
329 338
322 338
322 318
0 1 14 0 0 0 0 0 17 20 0 3
322 291
322 319
329 319
1 2 14 0 0 8320 0 4 13 0 0 3
214 337
214 291
488 291
0 1 16 0 0 4096 0 0 13 29 0 3
491 83
491 273
488 273
3 2 17 0 0 8320 0 18 16 0 0 4
385 243
469 243
469 93
520 93
0 2 18 0 0 8320 0 0 15 25 0 3
297 248
297 164
507 164
0 2 18 0 0 0 0 0 18 25 0 3
326 248
326 252
334 252
1 1 18 0 0 0 0 5 18 0 0 4
221 248
326 248
326 234
334 234
0 2 16 0 0 0 0 0 19 28 0 3
306 127
306 145
330 145
3 1 19 0 0 4224 0 19 15 0 0 4
381 136
504 136
504 155
507 155
0 1 16 0 0 0 0 0 19 29 0 3
306 83
306 127
330 127
1 1 16 0 0 8320 0 6 16 0 0 5
233 114
233 83
512 83
512 84
520 84
0
0
2049 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
2687728 1079360 100 100 0 0
0 0 0 0
1 66 162 136
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
12385 0
4 1 2
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
