CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 5 100 9
0 71 1280 680
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
16 C:\CM60S\BOM.DAT
0 7
0 71 1280 680
143654930 0
0
6 Title:
5 Name:
0
0
0
16
5 Lamp~
206 1156 72 0 2 3
11 9 2
0
0 0 624 0
3 100
-10 -24 11 -16
4 LAMP
-14 -22 14 -14
0
0
11 %D %1 %2 %V
0
0
0
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 L
8953 0 0
0
0
10 2-In NAND~
219 951 83 0 3 22
0 12 14 11
0
0 0 608 0
6 74LS00
-14 -24 28 -16
4 NAND
-7 -34 21 -26
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 2 0
1 U
4441 0 0
0
0
10 2-In NAND~
219 1031 86 0 3 22
0 11 10 9
0
0 0 608 0
6 74LS00
-14 -24 28 -16
4 NAND
-7 -34 21 -26
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 2 0
1 U
3618 0 0
0
0
10 2-In NAND~
219 947 150 0 3 22
0 14 13 12
0
0 0 608 0
6 74LS00
-14 -24 28 -16
4 NAND
-7 -33 21 -25
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 2 0
1 U
6153 0 0
0
0
10 2-In NAND~
219 1025 150 0 3 22
0 12 13 10
0
0 0 608 0
6 74LS00
-14 -24 28 -16
4 NAND
-7 -34 21 -26
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 2 0
1 U
5394 0 0
0
0
7 Ground~
168 1168 91 0 1 3
0 2
0
0 0 53344 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
7734 0 0
0
0
13 Logic Switch~
5 828 93 0 1 11
0 14
0
0 0 21344 0
2 0V
-7 -15 7 -7
2 V2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
9914 0 0
0
0
13 Logic Switch~
5 827 179 0 10 11
0 13 0 0 0 0 0 0 0 0
1
0
0 0 21344 0
2 5V
-7 -15 7 -7
2 V4
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
3747 0 0
0
0
13 Logic Switch~
5 288 298 0 10 11
0 3 0 0 0 0 0 0 0 0
1
0
0 0 21344 0
2 5V
-7 -15 7 -7
2 V1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3549 0 0
0
0
13 Logic Switch~
5 289 212 0 1 11
0 4
0
0 0 21344 0
2 0V
-7 -15 7 -7
2 V3
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
7931 0 0
0
0
10 2-In NAND~
219 343 238 0 3 22
0 4 3 5
0
0 0 608 0
6 74LS00
-14 -24 28 -16
4 NAND
-7 -33 21 -25
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 3 0
1 U
9325 0 0
0
0
10 2-In NAND~
219 393 321 0 3 22
0 5 3 6
0
0 0 608 0
6 74LS00
-14 -24 28 -16
4 NAND
-7 -34 21 -26
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 3 0
1 U
8903 0 0
0
0
10 2-In NAND~
219 607 254 0 3 22
0 7 6 8
0
0 0 608 0
6 74LS00
-14 -24 28 -16
4 NAND
-7 -34 21 -26
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 3 0
1 U
3834 0 0
0
0
10 2-In NAND~
219 400 168 0 3 22
0 4 5 7
0
0 0 608 0
6 74LS00
-14 -24 28 -16
4 NAND
-7 -34 21 -26
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 3 0
1 U
3363 0 0
0
0
7 Ground~
168 697 260 0 1 3
0 2
0
0 0 53344 0
0
4 GND2
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
7668 0 0
0
0
5 Lamp~
206 685 241 0 2 3
11 8 2
0
0 0 624 0
3 100
-10 -24 11 -16
4 LAMP
-14 -22 14 -14
0
0
11 %D %1 %2 %V
0
0
0
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 L
4718 0 0
0
0
20
3 1 9 0 0 16 0 3 1 0 0 3
1058 86
1058 85
1144 85
3 2 10 0 0 16 0 5 3 0 0 6
1052 150
1052 125
1009 125
1009 98
1007 98
1007 95
3 1 11 0 0 16 0 2 3 0 0 3
978 83
1007 83
1007 77
0 1 12 0 0 16 0 0 2 5 0 5
986 141
986 197
906 197
906 74
927 74
3 1 12 0 0 16 0 4 5 0 0 3
974 150
974 141
1001 141
0 2 13 0 0 16 0 0 5 9 0 3
923 179
1001 179
1001 159
0 2 14 0 0 16 0 0 2 8 0 3
887 93
887 92
927 92
1 1 14 0 0 16 0 7 4 0 0 4
840 93
887 93
887 141
923 141
1 2 13 0 0 16 0 8 4 0 0 3
839 179
923 179
923 159
1 2 2 0 0 16 0 6 1 0 0 2
1168 85
1168 85
1 2 3 0 0 4096 0 9 11 0 0 3
300 298
300 247
319 247
1 1 4 0 0 8192 0 10 11 0 0 3
301 212
301 229
319 229
0 2 5 0 0 4096 0 0 14 14 0 3
368 240
368 177
376 177
3 1 5 0 0 8320 0 11 12 0 0 4
370 238
368 238
368 312
369 312
1 2 3 0 0 8320 0 9 12 0 0 3
300 298
300 330
369 330
1 1 4 0 0 8320 0 10 14 0 0 3
301 212
301 159
376 159
3 2 6 0 0 4224 0 12 13 0 0 4
420 321
575 321
575 263
583 263
3 1 7 0 0 4224 0 14 13 0 0 4
427 168
575 168
575 245
583 245
3 1 8 0 0 4224 0 13 16 0 0 2
634 254
673 254
1 2 2 0 0 0 0 15 16 0 0 2
697 254
697 254
0
0
2049 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
788264 1079360 100 100 0 0
0 0 0 0
1 66 162 136
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
12385 0
4 2 2
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
