CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 9
32 88 1248 655
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
16 C:\CM60S\BOM.DAT
0 7
32 88 1248 655
143654930 0
0
6 Title:
5 Name:
0
0
0
17
13 Logic Switch~
5 191 311 0 1 11
0 5
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V4
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
8953 0 0
0
0
13 Logic Switch~
5 194 259 0 1 11
0 7
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V3
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
4441 0 0
0
0
13 Logic Switch~
5 191 203 0 1 11
0 9
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
3618 0 0
0
0
13 Logic Switch~
5 191 136 0 1 11
0 3
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
6153 0 0
0
0
7 Ground~
168 294 71 0 1 3
0 2
0
0 0 53360 180
0
4 GND5
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
5394 0 0
0
0
7 Ground~
168 521 317 0 1 3
0 2
0
0 0 53360 0
0
4 GND4
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
7734 0 0
0
0
7 Ground~
168 517 263 0 1 3
0 2
0
0 0 53360 0
0
4 GND3
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
9914 0 0
0
0
7 Ground~
168 518 210 0 1 3
0 2
0
0 0 53360 0
0
4 GND2
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
3747 0 0
0
0
7 Ground~
168 517 148 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
3549 0 0
0
0
9 2-In XOR~
219 343 309 0 3 22
0 6 5 4
0
0 0 624 0
6 74LS86
-21 -24 21 -16
3 U1D
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0
65 0 0 0 4 4 1 0
1 U
7931 0 0
0
0
9 2-In XOR~
219 344 254 0 3 22
0 8 7 6
0
0 0 624 0
6 74LS86
-21 -24 21 -16
3 U1C
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0
65 0 0 0 4 3 1 0
1 U
9325 0 0
0
0
9 2-In XOR~
219 343 201 0 3 22
0 10 9 8
0
0 0 624 0
6 74LS86
-21 -24 21 -16
3 U1B
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0
65 0 0 0 4 2 1 0
1 U
8903 0 0
0
0
9 2-In XOR~
219 341 143 0 3 22
0 2 3 10
0
0 0 624 0
6 74LS86
-21 -24 21 -16
3 U1A
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 389796381
65 0 0 0 4 1 1 0
1 U
3834 0 0
0
0
5 Lamp~
206 508 298 0 2 3
11 4 2
0
0 0 608 0
3 100
-10 -24 11 -16
2 L4
-7 -22 7 -14
0
0
11 %D %1 %2 %V
0
0
0
5

0 1 2 1 2 0
82 0 0 0 0 0 0 0
1 L
3363 0 0
0
0
5 Lamp~
206 505 244 0 2 3
11 6 2
0
0 0 608 0
3 100
-10 -24 11 -16
2 L3
-7 -22 7 -14
0
0
11 %D %1 %2 %V
0
0
0
5

0 1 2 1 2 0
82 0 0 0 0 0 0 0
1 L
7668 0 0
0
0
5 Lamp~
206 507 191 0 2 3
11 8 2
0
0 0 608 0
3 100
-10 -24 11 -16
2 L2
-7 -22 7 -14
0
0
11 %D %1 %2 %V
0
0
0
5

0 1 2 1 2 0
82 0 0 0 0 0 0 0
1 L
4718 0 0
0
0
5 Lamp~
206 507 130 0 2 3
11 10 2
0
0 0 608 0
3 100
-10 -24 11 -16
2 L1
-7 -22 7 -14
0
0
11 %D %1 %2 %V
0
0
0
5

0 1 2 1 2 0
82 0 0 0 0 0 0 0
1 L
3874 0 0
0
0
16
1 1 2 0 0 8320 0 13 5 0 0 3
325 134
294 134
294 79
1 2 3 0 0 8336 0 4 13 0 0 3
203 136
203 152
325 152
1 2 2 0 0 0 0 6 14 0 0 2
521 311
520 311
1 2 2 0 0 0 0 7 15 0 0 2
517 257
517 257
1 2 2 0 0 0 0 8 16 0 0 2
518 204
519 204
1 2 2 0 0 128 0 9 17 0 0 3
517 142
517 143
519 143
3 1 4 0 0 4224 0 10 14 0 0 4
376 309
488 309
488 311
496 311
1 2 5 0 0 4224 0 1 10 0 0 4
203 311
319 311
319 318
327 318
0 1 6 0 0 8192 0 0 10 10 0 5
396 254
396 280
319 280
319 300
327 300
3 1 6 0 0 4224 0 11 15 0 0 4
377 254
485 254
485 257
493 257
1 2 7 0 0 4224 0 2 11 0 0 4
206 259
320 259
320 263
328 263
0 1 8 0 0 8192 0 0 11 13 0 5
400 201
400 223
320 223
320 245
328 245
3 1 8 0 0 4224 0 12 16 0 0 4
376 201
487 201
487 204
495 204
1 2 9 0 0 8320 0 3 12 0 0 3
203 203
203 210
327 210
0 1 10 0 0 8192 0 0 12 16 0 5
403 143
403 171
319 171
319 192
327 192
3 1 10 0 0 4224 0 13 17 0 0 2
374 143
495 143
0
0
2049 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
3736738 1079360 100 100 0 0
0 0 0 0
1 66 162 136
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
12385 0
4 0.05 0.1
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
