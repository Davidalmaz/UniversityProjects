CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 10 1 100 9
2 87 647 629
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
16 C:\CM60S\BOM.DAT
0 7
2 87 647 629
143654930 0
0
6 Title:
5 Name:
0
0
0
19
13 Logic Switch~
5 123 293 0 10 11
0 3 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
4 CLK1
-12 -26 16 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
8953 0 0
0
0
13 Logic Switch~
5 30 92 0 1 11
0 6
0
0 0 21360 0
2 0V
-6 -16 8 -8
1 X
-3 -26 4 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
4441 0 0
0
0
7 Pulser~
4 54 316 0 10 12
0 16 17 18 19 0 0 5 5 2
7
0
0 0 4656 0
0
3 CLK
-10 -28 11 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
1 V
3618 0 0
0
0
2 +V
167 269 303 0 1 3
0 4
0
0 0 54256 512
2 5V
-7 -22 7 -14
2 V1
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
6153 0 0
0
0
9 2-In XOR~
219 444 159 0 3 22
0 5 9 8
0
0 0 624 0
6 74LS86
-21 -24 21 -16
3 U5B
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 4 0
1 U
5394 0 0
0
0
9 2-In XOR~
219 507 90 0 3 22
0 6 8 7
0
0 0 624 0
6 74LS86
-21 -24 21 -16
3 U5A
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 4 0
1 U
7734 0 0
0
0
7 Ground~
168 566 165 0 1 3
0 2
0
0 0 53360 0
0
4 GND4
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
9914 0 0
0
0
8 2-In OR~
219 186 205 0 3 22
0 13 12 11
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U4A
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 3 0
1 U
3747 0 0
0
0
9 Inverter~
13 84 190 0 2 22
0 6 14
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U3A
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 2 0
1 U
3549 0 0
0
0
9 2-In AND~
219 130 128 0 3 22
0 6 5 13
0
0 0 624 692
6 74LS08
-21 -24 21 -16
3 U2B
-14 -25 7 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 1 0
1 U
7931 0 0
0
0
9 2-In AND~
219 129 182 0 3 22
0 10 14 12
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U2A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 1 0
1 U
9325 0 0
0
0
7 Ground~
168 381 133 0 1 3
0 2
0
0 0 53360 0
0
4 GND3
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
8903 0 0
0
0
7 Ground~
168 390 204 0 1 3
0 2
0
0 0 53360 0
0
4 GND2
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3834 0 0
0
0
7 Ground~
168 197 103 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3363 0 0
0
0
6 74LS76
104 281 191 0 14 29
0 9 15 3 4 4 11 11 3 4
4 5 10 9 15
0
0 0 13040 0
6 74LS76
-21 -60 21 -52
2 U1
-7 -61 7 -53
0
15 DVCC=16;DGND=8;
131 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 4 16 1 2 3 9 12 6 7
8 15 14 11 10 4 16 1 2 3
9 12 6 7 8 15 14 11 10 0
65 0 0 0 1 0 0 0
1 U
7668 0 0
0
0
5 Lamp~
206 555 147 0 2 3
11 7 2
0
0 0 624 0
3 100
-10 -24 11 -16
1 Y
-4 -22 3 -14
0
0
11 %D %1 %2 %V
0
0
0
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 L
4718 0 0
0
0
5 Lamp~
206 369 114 0 2 3
11 5 2
0
0 0 624 0
3 100
-10 -24 11 -16
1 A
-4 -22 3 -14
0
0
11 %D %1 %2 %V
0
0
0
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 L
3874 0 0
0
0
5 Lamp~
206 378 186 0 2 3
11 9 2
0
0 0 624 0
3 100
-10 -24 11 -16
1 B
-4 -22 3 -14
0
0
11 %D %1 %2 %V
0
0
0
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 L
6671 0 0
0
0
5 Lamp~
206 185 87 0 2 3
11 6 2
0
0 0 624 0
3 100
-10 -24 11 -16
1 X
-4 -22 3 -14
0
0
11 %D %1 %2 %V
0
0
0
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 L
3789 0 0
0
0
30
8 0 3 0 0 4096 0 15 0 0 2 2
243 218
224 218
1 3 3 0 0 8320 0 1 15 0 0 4
135 293
224 293
224 173
243 173
10 0 4 0 0 4096 0 15 0 0 6 2
243 236
235 236
9 0 4 0 0 0 0 15 0 0 6 2
243 227
235 227
5 0 4 0 0 0 0 15 0 0 6 2
243 191
235 191
4 1 4 0 0 8320 0 15 4 0 0 5
243 182
235 182
235 320
269 320
269 312
1 0 5 0 0 4096 0 5 0 0 12 2
428 150
428 151
1 0 6 0 0 12416 0 6 0 0 15 5
491 81
492 81
492 32
76 32
76 100
3 1 7 0 0 8320 0 6 16 0 0 5
540 90
539 90
539 159
543 159
543 160
3 2 8 0 0 12416 0 5 6 0 0 5
477 159
477 158
476 158
476 99
491 99
2 0 9 0 0 28672 0 5 0 0 25 9
428 168
429 168
429 169
425 169
425 166
422 166
422 159
353 159
353 199
0 0 5 0 0 12288 0 0 0 28 0 5
350 153
351 153
351 151
428 151
428 148
0 2 5 0 0 8320 0 0 10 28 0 4
322 153
322 51
106 51
106 119
12 1 10 0 0 12432 0 15 11 0 0 6
319 164
325 164
325 252
102 252
102 173
105 173
1 0 6 0 0 0 0 19 0 0 17 2
173 100
61 100
1 0 6 0 0 0 0 10 0 0 17 2
106 137
61 137
1 1 6 0 0 0 0 2 9 0 0 4
42 92
61 92
61 190
69 190
0 7 11 0 0 8192 0 0 15 19 0 3
241 204
241 209
249 209
3 6 11 0 0 4224 0 8 15 0 0 5
219 205
235 205
235 204
249 204
249 200
3 2 12 0 0 8320 0 11 8 0 0 4
150 182
156 182
156 214
173 214
3 1 13 0 0 8320 0 10 8 0 0 4
151 128
165 128
165 196
173 196
2 2 14 0 0 4224 0 9 11 0 0 2
105 190
105 191
14 2 15 0 0 8320 0 15 15 0 0 6
319 209
330 209
330 88
230 88
230 164
249 164
0 1 9 0 0 4224 0 0 15 25 0 4
340 199
340 65
249 65
249 155
13 1 9 0 0 0 0 15 18 0 0 3
313 200
313 199
366 199
1 2 2 0 0 4096 0 7 16 0 0 4
566 159
568 159
568 160
567 160
1 2 2 0 0 0 0 12 17 0 0 2
381 127
381 127
11 1 5 0 0 0 0 15 17 0 0 5
313 155
313 153
350 153
350 127
357 127
1 2 2 0 0 0 0 13 18 0 0 2
390 198
390 199
1 2 2 0 0 4224 0 14 19 0 0 2
197 97
197 100
0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
