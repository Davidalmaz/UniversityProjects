CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 9
7 78 1223 645
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
16 C:\CM60S\BOM.DAT
0 7
7 78 1223 645
143654930 0
0
6 Title:
5 Name:
0
0
0
32
7 Ground~
168 781 369 0 1 3
0 0
0
0 0 53344 0
0
4 GND4
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
8953 0 0
0
0
13 Logic Switch~
5 279 317 0 1 11
0 17
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 Z1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
4441 0 0
0
0
13 Logic Switch~
5 41 210 0 1 11
0 15
0
0 0 21360 0
2 0V
-6 -16 8 -8
1 Z
-3 -26 4 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3618 0 0
0
0
13 Logic Switch~
5 37 68 0 1 11
0 22
0
0 0 21360 0
2 0V
-6 -16 8 -8
1 X
-3 -26 4 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
6153 0 0
0
0
13 Logic Switch~
5 42 151 0 1 11
0 21
0
0 0 21360 0
2 0V
-10 -16 4 -8
1 Y
-3 -26 4 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5394 0 0
0
0
13 Logic Switch~
5 241 405 0 1 11
0 18
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 X1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
7734 0 0
0
0
13 Logic Switch~
5 247 361 0 1 11
0 16
0
0 0 21360 0
2 0V
-10 -16 4 -8
2 Y1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
9914 0 0
0
0
10 3-In NAND~
219 724 361 0 4 22
0 3 13 12 14
0
0 0 624 0
6 74LS10
-21 -28 21 -20
3 U8C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
17

0 9 10 11 8 1 2 13 12 3
4 5 6 9 10 11 8 0
65 0 0 0 3 3 7 0
1 U
3747 0 0
0
0
10 3-In NAND~
219 557 452 0 4 22
0 6 5 4 12
0
0 0 624 0
6 74LS10
-21 -28 21 -20
3 U8B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
17

0 3 4 5 6 1 2 13 12 3
4 5 6 9 10 11 8 0
65 0 0 0 3 2 7 0
1 U
3549 0 0
0
0
10 3-In NAND~
219 647 374 0 4 22
0 9 8 7 13
0
0 0 624 0
6 74LS10
-21 -28 21 -20
3 U8A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
17

0 1 2 13 12 1 2 13 12 3
4 5 6 9 10 11 8 0
65 0 0 0 3 1 7 0
1 U
7931 0 0
0
0
10 3-In NAND~
219 554 298 0 4 22
0 11 10 4 3
0
0 0 624 0
6 74LS10
-21 -28 21 -20
3 U6C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
17

0 9 10 11 8 1 2 13 12 3
4 5 6 9 10 11 8 0
65 0 0 0 3 3 5 0
1 U
9325 0 0
0
0
7 Ground~
168 367 422 0 1 3
0 2
0
0 0 53360 0
0
4 GND5
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
8903 0 0
0
0
7 Ground~
168 1057 200 0 1 3
0 2
0
0 0 53360 0
0
4 GND3
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3834 0 0
0
0
10 2-In NAND~
219 903 118 0 3 22
0 22 21 24
0
0 0 624 0
6 74LS00
-14 -24 28 -16
3 U5A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 4 0
1 U
3363 0 0
0
0
10 3-In NAND~
219 893 234 0 4 22
0 19 20 15 23
0
0 0 624 0
6 74LS10
-21 -28 21 -20
3 U3C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
17

0 9 10 11 8 1 2 13 12 3
4 5 6 9 10 11 8 0
65 0 0 0 3 3 2 0
1 U
7668 0 0
0
0
10 2-In NAND~
219 1003 192 0 3 22
0 24 23 25
0
0 0 624 0
6 74LS00
-14 -24 28 -16
3 U5B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 4 0
1 U
4718 0 0
0
0
10 2-In NAND~
219 596 89 0 3 22
0 19 21 28
0
0 0 624 0
6 74LS00
-14 -24 28 -16
3 U4D
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 3 0
1 U
3874 0 0
0
0
7 Ground~
168 749 178 0 1 3
0 2
0
0 0 53360 0
0
4 GND2
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
6671 0 0
0
0
10 3-In NAND~
219 588 213 0 4 22
0 22 20 26 27
0
0 0 624 0
6 74LS10
-21 -28 21 -20
3 U3B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
17

0 3 4 5 6 1 2 13 12 3
4 5 6 9 10 11 8 0
65 0 0 0 3 2 2 0
1 U
3789 0 0
0
0
10 2-In NAND~
219 698 171 0 3 22
0 28 27 29
0
0 0 624 0
6 74LS00
-14 -24 28 -16
3 U4C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 3 0
1 U
4871 0 0
0
0
7 Ground~
168 485 163 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3750 0 0
0
0
10 2-In NAND~
219 438 158 0 3 22
0 32 31 30
0
0 0 624 0
6 74LS00
-14 -24 28 -16
3 U4A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 3 0
1 U
8778 0 0
0
0
10 2-In NAND~
219 312 114 0 3 22
0 22 15 32
0
0 0 624 0
6 74LS00
-14 -24 28 -16
3 U2D
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 1 0
1 U
538 0 0
0
0
10 2-In NAND~
219 245 154 0 3 22
0 21 21 20
0
0 0 624 0
6 74LS00
-14 -24 28 -16
3 U2C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 1 0
1 U
6843 0 0
0
0
10 2-In NAND~
219 248 244 0 3 22
0 15 15 26
0
0 0 624 0
6 74LS00
-14 -24 28 -16
3 U2B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 1 0
1 U
3136 0 0
0
0
10 3-In NAND~
219 366 196 0 4 22
0 19 20 26 31
0
0 0 624 0
6 74LS10
-21 -28 21 -20
3 U3A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
17

0 1 2 13 12 1 2 13 12 3
4 5 6 9 10 11 8 0
65 0 0 0 3 1 2 0
1 U
5950 0 0
0
0
10 2-In NAND~
219 258 62 0 3 22
0 22 22 19
0
0 0 624 0
6 74LS00
-14 -24 28 -16
3 U2A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 1 0
1 U
5670 0 0
0
0
7 74LS155
120 406 355 0 14 29
0 17 17 16 18 2 2 11 6 9
8 7 10 5 4
0
0 0 13040 0
7 74LS155
-24 -51 25 -43
2 U1
-7 -52 7 -44
0
15 DVCC=16;DGND=8;
114 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 2 3 13 14 15 4 5 6
7 12 11 10 9 1 2 3 13 14
15 4 5 6 7 12 11 10 9 0
65 0 0 0 1 0 0 0
1 U
6828 0 0
0
0
5 Lamp~
206 771 350 0 2 3
11 14 2
0
0 0 624 0
3 100
-10 -24 11 -16
2 L5
-7 -22 7 -14
0
0
11 %D %1 %2 %V
0
0
0
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 L
6735 0 0
0
0
5 Lamp~
206 1047 181 0 2 3
11 25 2
0
0 0 624 0
3 100
-10 -24 11 -16
2 L3
-7 -22 7 -14
0
0
11 %D %1 %2 %V
0
0
0
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 L
8365 0 0
0
0
5 Lamp~
206 739 159 0 2 3
11 29 2
0
0 0 624 0
3 100
-10 -24 11 -16
2 L2
-7 -22 7 -14
0
0
11 %D %1 %2 %V
0
0
0
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 L
4132 0 0
0
0
5 Lamp~
206 475 144 0 2 3
11 30 2
0
0 0 624 0
3 100
-10 -24 11 -16
2 L1
-7 -22 7 -14
0
0
11 %D %1 %2 %V
0
0
0
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 L
4551 0 0
0
0
55
1 2 0 0 0 0 0 1 29 0 0 2
781 363
783 363
0 3 4 0 0 4112 0 0 9 8 0 3
472 391
472 461
533 461
13 2 5 0 0 8320 0 28 9 0 0 4
444 382
486 382
486 452
533 452
8 1 6 0 0 8320 0 28 9 0 0 4
444 337
503 337
503 443
533 443
11 3 7 0 0 4224 0 28 10 0 0 4
444 364
492 364
492 383
623 383
10 2 8 0 0 4224 0 28 10 0 0 4
444 355
492 355
492 374
623 374
9 1 9 0 0 4224 0 28 10 0 0 4
444 346
492 346
492 365
623 365
14 3 4 0 0 8320 0 28 11 0 0 4
444 391
520 391
520 307
530 307
12 2 10 0 0 8320 0 28 11 0 0 4
444 373
507 373
507 298
530 298
7 1 11 0 0 4224 0 28 11 0 0 4
444 328
494 328
494 289
530 289
4 3 12 0 0 4224 0 9 8 0 0 4
584 452
695 452
695 370
700 370
4 2 13 0 0 4224 0 10 8 0 0 4
674 374
676 374
676 361
700 361
4 1 3 0 0 128 0 11 8 0 0 4
581 298
571 298
571 352
700 352
1 4 14 0 0 8320 0 29 8 0 0 3
759 363
759 361
751 361
0 1 15 0 0 8192 0 0 3 50 0 3
218 215
218 210
53 210
1 0 16 0 0 0 0 7 0 0 20 2
259 361
259 361
1 0 2 0 0 0 0 12 0 0 18 3
367 416
368 415
368 391
5 6 2 0 0 4224 0 28 28 0 0 2
368 382
368 391
1 0 17 0 0 16512 0 2 0 0 22 7
291 317
291 316
290 316
290 318
363 318
363 333
368 333
0 3 16 0 0 4224 0 0 28 0 0 4
255 361
360 361
360 355
374 355
1 4 18 0 0 12416 0 6 28 0 0 6
253 405
255 405
255 403
360 403
360 364
374 364
1 2 17 0 0 128 0 28 28 0 0 3
374 328
368 328
368 337
0 1 19 0 0 4224 0 0 15 39 0 4
344 62
861 62
861 225
869 225
0 2 20 0 0 8320 0 0 15 34 0 3
533 216
533 234
869 234
2 3 15 0 0 20608 0 23 15 0 0 7
288 123
284 123
284 215
281 215
281 272
869 272
869 243
0 2 21 0 0 8192 0 0 14 38 0 3
554 94
554 127
879 127
0 1 22 0 0 8320 0 0 14 35 0 3
532 204
532 109
879 109
4 2 23 0 0 4224 0 15 16 0 0 4
920 234
971 234
971 201
979 201
3 1 24 0 0 8320 0 14 16 0 0 4
930 118
971 118
971 183
979 183
1 3 25 0 0 4224 0 0 16 32 0 3
1035 194
1030 194
1030 192
1 2 2 0 0 128 0 13 30 0 0 2
1057 194
1059 194
1 3 25 0 0 0 0 30 0 0 30 4
1035 194
1035 195
1033 195
1033 194
0 3 26 0 0 4224 0 0 19 44 0 3
332 244
564 244
564 222
0 2 20 0 0 0 0 0 19 45 0 5
304 154
304 216
556 216
556 213
564 213
0 1 22 0 0 0 0 0 19 55 0 5
273 105
273 144
459 144
459 204
564 204
4 2 27 0 0 4224 0 19 20 0 0 4
615 213
666 213
666 180
674 180
3 1 28 0 0 8320 0 17 20 0 0 4
623 89
666 89
666 162
674 162
0 2 21 0 0 12416 0 0 17 51 0 6
214 144
217 144
217 94
564 94
564 98
572 98
0 1 19 0 0 0 0 0 17 46 0 3
344 62
344 80
572 80
1 2 2 0 0 0 0 18 31 0 0 2
749 172
751 172
1 3 29 0 0 8320 0 31 20 0 0 4
727 172
727 173
725 173
725 171
1 2 2 0 0 0 0 21 32 0 0 2
485 157
487 157
1 3 30 0 0 8320 0 32 22 0 0 3
463 157
463 158
465 158
3 3 26 0 0 0 0 25 26 0 0 4
275 244
334 244
334 205
342 205
3 2 20 0 0 0 0 24 26 0 0 4
272 154
334 154
334 196
342 196
3 1 19 0 0 0 0 27 26 0 0 4
285 62
344 62
344 187
342 187
4 2 31 0 0 4224 0 26 22 0 0 3
393 196
393 167
414 167
3 1 32 0 0 4224 0 23 22 0 0 4
339 114
393 114
393 149
414 149
2 0 15 0 0 0 0 25 0 0 50 6
224 253
225 253
225 253
217 253
217 235
218 235
0 1 15 0 0 0 0 0 25 25 0 4
281 215
218 215
218 235
224 235
0 1 21 0 0 0 0 0 24 52 0 3
214 164
214 144
222 144
1 2 21 0 0 0 0 5 24 0 0 8
54 151
63 151
63 163
97 163
97 164
214 164
214 163
221 163
0 2 22 0 0 0 0 0 27 54 0 3
225 72
225 71
234 71
0 1 22 0 0 0 0 0 27 55 0 3
225 105
225 53
234 53
1 1 22 0 0 0 0 4 23 0 0 6
49 68
58 68
58 106
225 106
225 105
288 105
0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
