CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 570 30 100 9
32 88 1248 655
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
16 C:\CM60S\BOM.DAT
0 7
32 88 1248 655
143654930 0
0
6 Title:
5 Name:
0
0
0
48
13 Logic Switch~
5 310 766 0 1 11
0 5
0
0 0 21360 0
2 0V
-6 -16 8 -8
3 V15
-9 -26 12 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
8953 0 0
0
0
13 Logic Switch~
5 309 816 0 1 11
0 5
0
0 0 21360 0
2 0V
-6 -16 8 -8
3 V14
-9 -26 12 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
4441 0 0
0
0
13 Logic Switch~
5 309 863 0 1 11
0 5
0
0 0 21360 0
2 0V
-6 -16 8 -8
3 V13
-9 -26 12 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
3618 0 0
0
0
13 Logic Switch~
5 311 907 0 1 11
0 5
0
0 0 21360 0
2 0V
-6 -16 8 -8
3 V12
-9 -26 12 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
6153 0 0
0
0
13 Logic Switch~
5 310 949 0 1 11
0 5
0
0 0 21360 0
2 0V
-6 -16 8 -8
3 V11
-9 -26 12 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
5394 0 0
0
0
13 Logic Switch~
5 827 291 0 1 11
0 13
0
0 0 21360 0
2 0V
-6 -16 8 -8
3 V10
-9 -26 12 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
7734 0 0
0
0
13 Logic Switch~
5 826 341 0 1 11
0 13
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V9
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
9914 0 0
0
0
13 Logic Switch~
5 826 388 0 1 11
0 13
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V8
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
3747 0 0
0
0
13 Logic Switch~
5 828 432 0 1 11
0 13
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V7
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
3549 0 0
0
0
13 Logic Switch~
5 827 474 0 1 11
0 13
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V6
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
7931 0 0
0
0
13 Logic Switch~
5 310 476 0 1 11
0 19
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V5
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
9325 0 0
0
0
13 Logic Switch~
5 311 434 0 1 11
0 19
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V4
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
8903 0 0
0
0
13 Logic Switch~
5 309 390 0 1 11
0 19
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V3
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
3834 0 0
0
0
13 Logic Switch~
5 309 343 0 1 11
0 19
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
3363 0 0
0
0
13 Logic Switch~
5 310 293 0 1 11
0 19
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
7668 0 0
0
0
6 74LS83
105 437 626 0 14 29
0 2 4 2 2 3 2 2 3 5
10 9 8 7 6
0
0 0 13040 0
7 74LS83A
-24 -60 25 -52
2 U3
-7 -61 7 -53
0
15 DVCC=5;DGND=12;
125 %D [%5bi %12bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 3 8 10 16 4 7 11 13
15 2 6 9 14 1 3 8 10 16
4 7 11 13 15 2 6 9 14 0
65 0 0 0 1 0 0 0
1 U
4718 0 0
0
0
7 Ground~
168 641 652 0 1 3
0 2
0
0 0 53360 90
0
4 GND9
-14 -28 14 -20
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
3874 0 0
0
0
9 V Source~
197 274 577 0 2 5
0 4 2
0
0 0 17264 0
3 10V
13 0 34 8
3 Vs6
13 -10 34 -2
0
0
11 %D %1 %2 %V
0
0
0
5

0 1 2 1 2 0
86 0 0 0 0 0 0 0
2 Vs
6671 0 0
0
0
7 Ground~
168 328 607 0 1 3
0 2
0
0 0 53360 0
0
4 GND8
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
3789 0 0
0
0
9 V Source~
197 284 662 0 2 5
0 3 2
0
0 0 17264 0
3 10V
13 0 34 8
3 Vs5
13 -10 34 -2
0
0
11 %D %1 %2 %V
0
0
0
5

0 1 2 1 2 0
86 0 0 0 0 0 0 0
2 Vs
4871 0 0
0
0
7 Ground~
168 339 695 0 1 3
0 2
0
0 0 53360 0
0
4 GND7
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
3750 0 0
0
0
6 74LS83
105 954 151 0 14 29
0 12 12 2 2 11 11 2 2 13
18 17 16 15 14
0
0 0 13040 0
7 74LS83A
-24 -60 25 -52
2 U2
-7 -61 7 -53
0
15 DVCC=5;DGND=12;
125 %D [%5bi %12bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 3 8 10 16 4 7 11 13
15 2 6 9 14 1 3 8 10 16
4 7 11 13 15 2 6 9 14 0
65 0 0 0 1 0 0 0
1 U
8778 0 0
0
0
7 Ground~
168 1158 177 0 1 3
0 2
0
0 0 53360 90
0
4 GND6
-14 -28 14 -20
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
538 0 0
0
0
9 V Source~
197 791 102 0 2 5
0 12 2
0
0 0 17264 0
3 10V
13 0 34 8
3 Vs4
13 -10 34 -2
0
0
11 %D %1 %2 %V
0
0
0
5

0 1 2 1 2 0
86 0 0 0 0 0 0 0
2 Vs
6843 0 0
0
0
7 Ground~
168 845 132 0 1 3
0 2
0
0 0 53360 0
0
4 GND5
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
3136 0 0
0
0
9 V Source~
197 801 187 0 2 5
0 11 2
0
0 0 17264 0
3 10V
13 0 34 8
3 Vs3
13 -10 34 -2
0
0
11 %D %1 %2 %V
0
0
0
5

0 1 2 1 2 0
86 0 0 0 0 0 0 0
2 Vs
5950 0 0
0
0
7 Ground~
168 856 220 0 1 3
0 2
0
0 0 53360 0
0
4 GND4
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
5670 0 0
0
0
7 Ground~
168 339 222 0 1 3
0 2
0
0 0 53360 0
0
4 GND3
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
6828 0 0
0
0
9 V Source~
197 284 189 0 2 5
0 20 2
0
0 0 17264 0
3 10V
13 0 34 8
3 Vs2
13 -10 34 -2
0
0
11 %D %1 %2 %V
0
0
0
5

0 1 2 1 2 0
86 0 0 0 0 0 0 0
2 Vs
6735 0 0
0
0
7 Ground~
168 328 134 0 1 3
0 2
0
0 0 53360 0
0
4 GND2
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
8365 0 0
0
0
9 V Source~
197 274 104 0 2 5
0 21 2
0
0 0 17264 0
3 10V
13 0 34 8
3 Vs1
13 -10 34 -2
0
0
11 %D %1 %2 %V
0
0
0
5

0 1 2 1 2 0
86 0 0 0 0 0 0 0
2 Vs
4132 0 0
0
0
7 Ground~
168 641 179 0 1 3
0 2
0
0 0 53360 90
0
4 GND1
-14 -28 14 -20
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
4551 0 0
0
0
6 74LS83
105 437 153 0 14 29
0 2 21 2 21 20 20 2 2 19
26 25 24 23 22
0
0 0 13040 0
7 74LS83A
-24 -60 25 -52
2 U1
-7 -61 7 -53
0
15 DVCC=5;DGND=12;
125 %D [%5bi %12bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 3 8 10 16 4 7 11 13
15 2 6 9 14 1 3 8 10 16
4 7 11 13 15 2 6 9 14 0
65 0 0 0 1 0 0 0
1 U
3635 0 0
0
0
5 Lamp~
206 549 562 0 2 3
11 10 2
0
0 0 608 0
3 100
-10 -24 11 -16
2 s8
-7 -22 7 -14
0
0
11 %D %1 %2 %V
0
0
0
5

0 1 2 1 2 0
82 0 0 0 0 0 0 0
1 L
3973 0 0
0
0
5 Lamp~
206 550 602 0 2 3
11 9 2
0
0 0 608 0
3 100
-10 -24 11 -16
2 s7
-7 -22 7 -14
0
0
11 %D %1 %2 %V
0
0
0
5

0 1 2 1 2 0
82 0 0 0 0 0 0 0
1 L
3851 0 0
0
0
5 Lamp~
206 551 641 0 2 3
11 8 2
0
0 0 608 0
3 100
-10 -24 11 -16
2 s6
-7 -22 7 -14
0
0
11 %D %1 %2 %V
0
0
0
5

0 1 2 1 2 0
82 0 0 0 0 0 0 0
1 L
8383 0 0
0
0
5 Lamp~
206 551 681 0 2 3
11 7 2
0
0 0 608 0
3 100
-10 -24 11 -16
2 s5
-7 -22 7 -14
0
0
11 %D %1 %2 %V
0
0
0
5

0 1 2 1 2 0
82 0 0 0 0 0 0 0
1 L
9334 0 0
0
0
5 Lamp~
206 550 515 0 2 3
11 6 2
0
0 0 608 0
3 100
-10 -24 11 -16
7 ACARREO
-24 -22 25 -14
0
0
11 %D %1 %2 %V
0
0
0
5

0 1 2 1 2 0
82 0 0 0 0 0 0 0
1 L
7471 0 0
0
0
5 Lamp~
206 1066 87 0 2 3
11 18 2
0
0 0 608 0
3 100
-10 -24 11 -16
2 s4
-7 -22 7 -14
0
0
11 %D %1 %2 %V
0
0
0
5

0 1 2 1 2 0
82 0 0 0 0 0 0 0
1 L
3334 0 0
0
0
5 Lamp~
206 1067 127 0 2 3
11 17 2
0
0 0 608 0
3 100
-10 -24 11 -16
2 s3
-7 -22 7 -14
0
0
11 %D %1 %2 %V
0
0
0
5

0 1 2 1 2 0
82 0 0 0 0 0 0 0
1 L
3559 0 0
0
0
5 Lamp~
206 1068 166 0 2 3
11 16 2
0
0 0 608 0
3 100
-10 -24 11 -16
2 s2
-7 -22 7 -14
0
0
11 %D %1 %2 %V
0
0
0
5

0 1 2 1 2 0
82 0 0 0 0 0 0 0
1 L
984 0 0
0
0
5 Lamp~
206 1068 206 0 2 3
11 15 2
0
0 0 608 0
3 100
-10 -24 11 -16
2 s1
-7 -22 7 -14
0
0
11 %D %1 %2 %V
0
0
0
5

0 1 2 1 2 0
82 0 0 0 0 0 0 0
1 L
7557 0 0
0
0
5 Lamp~
206 1067 36 0 2 3
11 14 2
0
0 0 608 0
3 100
-10 -24 11 -16
7 ACARREO
-24 -22 25 -14
0
0
11 %D %1 %2 %V
0
0
0
5

0 1 2 1 2 0
82 0 0 0 0 0 0 0
1 L
3146 0 0
0
0
5 Lamp~
206 550 42 0 2 3
11 22 2
0
0 0 608 0
3 100
-10 -24 11 -16
7 ACARREO
-24 -22 25 -14
0
0
11 %D %1 %2 %V
0
0
0
5

0 1 2 1 2 0
82 0 0 0 0 0 0 0
1 L
5687 0 0
0
0
5 Lamp~
206 551 208 0 2 3
11 23 2
0
0 0 608 0
3 100
-10 -24 11 -16
2 s1
-7 -22 7 -14
0
0
11 %D %1 %2 %V
0
0
0
5

0 1 2 1 2 0
82 0 0 0 0 0 0 0
1 L
7939 0 0
0
0
5 Lamp~
206 551 168 0 2 3
11 24 2
0
0 0 608 0
3 100
-10 -24 11 -16
2 s2
-7 -22 7 -14
0
0
11 %D %1 %2 %V
0
0
0
5

0 1 2 1 2 0
82 0 0 0 0 0 0 0
1 L
3308 0 0
0
0
5 Lamp~
206 550 129 0 2 3
11 25 2
0
0 0 608 0
3 100
-10 -24 11 -16
2 s3
-7 -22 7 -14
0
0
11 %D %1 %2 %V
0
0
0
5

0 1 2 1 2 0
82 0 0 0 0 0 0 0
1 L
3408 0 0
0
0
5 Lamp~
206 549 89 0 2 3
11 26 2
0
0 0 608 0
3 100
-10 -24 11 -16
2 s4
-7 -22 7 -14
0
0
11 %D %1 %2 %V
0
0
0
5

0 1 2 1 2 0
82 0 0 0 0 0 0 0
1 L
9773 0 0
0
0
75
0 5 3 0 0 8192 0 0 16 2 0 3
373 637
373 626
405 626
1 8 3 0 0 8320 0 20 16 0 0 5
284 641
284 637
397 637
397 653
405 653
0 6 2 0 0 8192 0 0 16 4 0 3
393 644
393 635
405 635
1 7 2 0 0 8192 0 21 16 0 0 3
339 689
339 644
405 644
1 2 4 0 0 8320 0 18 16 0 0 5
274 556
274 552
397 552
397 599
405 599
0 1 2 0 0 0 0 0 16 8 0 3
395 597
395 590
405 590
0 3 2 0 0 0 0 0 16 8 0 3
397 607
397 608
405 608
0 4 2 0 0 8192 0 0 16 15 0 5
326 596
326 597
397 597
397 617
405 617
1 0 5 0 0 4096 0 5 0 0 10 3
322 949
397 949
397 907
1 0 5 0 0 0 0 4 0 0 11 3
323 907
397 907
397 863
1 0 5 0 0 4096 0 3 0 0 12 3
321 863
397 863
397 816
1 0 5 0 0 0 0 2 0 0 13 3
321 816
397 816
397 766
1 9 5 0 0 8320 0 1 16 0 0 4
322 766
397 766
397 671
405 671
2 1 2 0 0 16 0 20 21 0 0 6
284 683
284 688
326 688
326 685
339 685
339 689
2 1 2 0 0 0 0 18 19 0 0 6
274 598
274 603
315 603
315 596
328 596
328 601
2 0 2 0 0 0 0 37 0 0 18 3
563 694
602 694
602 654
2 0 2 0 0 8192 0 38 0 0 19 4
562 528
624 528
624 653
629 653
2 0 2 0 0 0 0 35 0 0 20 3
562 615
602 615
602 654
2 0 2 0 0 0 0 34 0 0 20 3
561 575
629 575
629 653
2 1 2 0 0 0 0 36 17 0 0 4
563 654
626 654
626 653
634 653
14 1 6 0 0 4224 0 16 38 0 0 3
469 671
469 528
538 528
13 1 7 0 0 8320 0 16 37 0 0 4
469 644
504 644
504 694
539 694
12 1 8 0 0 4224 0 16 36 0 0 4
469 635
531 635
531 654
539 654
11 1 9 0 0 4224 0 16 35 0 0 4
469 626
530 626
530 615
538 615
10 1 10 0 0 8320 0 16 34 0 0 3
469 617
469 575
537 575
0 8 2 0 0 0 0 0 22 27 0 3
908 169
908 178
922 178
0 7 2 0 0 0 0 0 22 39 0 3
856 209
856 169
922 169
0 6 11 0 0 8192 0 0 22 29 0 3
896 151
896 160
922 160
1 5 11 0 0 8320 0 26 22 0 0 3
801 166
801 151
922 151
0 4 2 0 0 0 0 0 22 31 0 4
883 133
914 133
914 142
922 142
0 3 2 0 0 0 0 0 22 40 0 5
845 121
845 119
883 119
883 133
922 133
0 2 12 0 0 4096 0 0 22 33 0 3
892 77
892 124
922 124
1 1 12 0 0 8320 0 24 22 0 0 5
791 81
791 77
914 77
914 115
922 115
1 0 13 0 0 4096 0 10 0 0 35 3
839 474
914 474
914 432
1 0 13 0 0 0 0 9 0 0 36 3
840 432
914 432
914 388
1 0 13 0 0 4096 0 8 0 0 37 3
838 388
914 388
914 341
1 0 13 0 0 0 0 7 0 0 38 3
838 341
914 341
914 291
1 9 13 0 0 8320 0 6 22 0 0 4
839 291
914 291
914 196
922 196
2 1 2 0 0 0 0 26 27 0 0 6
801 208
801 213
843 213
843 209
856 209
856 214
2 1 2 0 0 0 0 24 25 0 0 6
791 123
791 128
832 128
832 121
845 121
845 126
2 0 2 0 0 0 0 42 0 0 43 3
1080 219
1119 219
1119 179
2 0 2 0 0 8320 0 43 0 0 44 4
1079 49
1141 49
1141 178
1146 178
2 0 2 0 0 0 0 40 0 0 45 3
1079 140
1119 140
1119 179
2 0 2 0 0 0 0 39 0 0 45 3
1078 100
1146 100
1146 178
2 1 2 0 0 0 0 41 23 0 0 4
1080 179
1143 179
1143 178
1151 178
14 1 14 0 0 4224 0 22 43 0 0 3
986 196
986 49
1055 49
13 1 15 0 0 8320 0 22 42 0 0 4
986 169
1021 169
1021 219
1056 219
12 1 16 0 0 4224 0 22 41 0 0 4
986 160
1048 160
1048 179
1056 179
11 1 17 0 0 4224 0 22 40 0 0 4
986 151
1047 151
1047 140
1055 140
10 1 18 0 0 8320 0 22 39 0 0 3
986 142
986 100
1054 100
1 0 19 0 0 4096 0 11 0 0 52 3
322 476
397 476
397 434
1 0 19 0 0 0 0 12 0 0 53 3
323 434
397 434
397 390
1 0 19 0 0 4096 0 13 0 0 54 3
321 390
397 390
397 343
1 0 19 0 0 0 0 14 0 0 55 3
321 343
397 343
397 293
1 9 19 0 0 8320 0 15 33 0 0 4
322 293
397 293
397 198
405 198
0 7 2 0 0 0 0 0 33 57 0 3
376 180
376 171
405 171
0 8 2 0 0 0 0 0 33 64 0 3
339 211
339 180
405 180
0 6 20 0 0 8192 0 0 33 59 0 3
392 153
392 162
405 162
1 5 20 0 0 8320 0 29 33 0 0 3
284 168
284 153
405 153
0 1 2 0 0 0 0 0 33 61 0 4
376 109
376 88
405 88
405 117
0 3 2 0 0 0 0 0 33 65 0 5
326 123
326 109
397 109
397 135
405 135
0 2 21 0 0 4096 0 0 33 63 0 4
360 123
397 123
397 126
405 126
1 4 21 0 0 8320 0 31 33 0 0 5
274 83
274 79
360 79
360 144
405 144
2 1 2 0 0 0 0 29 28 0 0 6
284 210
284 215
326 215
326 211
339 211
339 216
2 1 2 0 0 0 0 31 30 0 0 6
274 125
274 130
315 130
315 123
328 123
328 128
2 0 2 0 0 0 0 45 0 0 68 3
563 221
602 221
602 181
2 0 2 0 0 128 0 44 0 0 69 4
562 55
624 55
624 180
629 180
2 0 2 0 0 0 0 47 0 0 70 3
562 142
602 142
602 181
2 0 2 0 0 0 0 48 0 0 70 3
561 102
629 102
629 180
2 1 2 0 0 0 0 46 32 0 0 4
563 181
626 181
626 180
634 180
14 1 22 0 0 4224 0 33 44 0 0 3
469 198
469 55
538 55
13 1 23 0 0 8320 0 33 45 0 0 4
469 171
504 171
504 221
539 221
12 1 24 0 0 4224 0 33 46 0 0 4
469 162
531 162
531 181
539 181
11 1 25 0 0 4224 0 33 47 0 0 4
469 153
530 153
530 142
538 142
10 1 26 0 0 8320 0 33 48 0 0 3
469 144
469 102
537 102
6
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 4
226 646 266 670
236 654 268 670
4 1001
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 4
212 561 252 585
222 569 254 585
4 0100
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 4
735 91 775 115
745 99 777 115
4 1100
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 4
744 171 784 195
754 179 786 195
4 1100
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 4
227 173 267 197
237 181 269 197
4 1100
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 4
220 89 260 113
230 97 262 113
4 0101
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
