CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 9
0 71 1280 672
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
16 C:\CM60S\BOM.DAT
0 7
0 71 1280 672
143654930 0
0
6 Title:
5 Name:
0
0
0
28
13 Logic Switch~
5 89 336 0 10 11
0 27 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V5
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
8953 0 0
0
0
13 Logic Switch~
5 72 294 0 1 11
0 19
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V4
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
4441 0 0
0
0
13 Logic Switch~
5 70 244 0 1 11
0 20
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V3
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3618 0 0
0
0
13 Logic Switch~
5 67 186 0 1 11
0 21
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
6153 0 0
0
0
13 Logic Switch~
5 66 129 0 10 11
0 22 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5394 0 0
0
0
9 Inverter~
13 577 159 0 2 22
0 5 4
0
0 0 624 782
6 74LS04
-21 -19 21 -11
3 U5D
16 -8 37 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 9 8 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 4 4 0
1 U
7734 0 0
0
0
9 2-In AND~
219 497 155 0 3 22
0 8 7 11
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U1D
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 1 0
1 U
9914 0 0
0
0
9 2-In AND~
219 494 78 0 3 22
0 10 9 12
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U6A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 5 0
1 U
3747 0 0
0
0
9 2-In AND~
219 547 112 0 3 22
0 12 11 5
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U6B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 5 0
1 U
3549 0 0
0
0
7 Ground~
168 803 197 0 1 3
0 2
0
0 0 53360 0
0
4 GND7
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
7931 0 0
0
0
9 2-In XOR~
219 186 263 0 3 22
0 19 27 23
0
0 0 624 0
6 74LS86
-21 -24 21 -16
3 U3A
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 3 0
1 U
9325 0 0
0
0
9 2-In XOR~
219 189 221 0 3 22
0 20 27 24
0
0 0 624 0
6 74LS86
-21 -24 21 -16
3 U3B
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 3 0
1 U
8903 0 0
0
0
9 2-In XOR~
219 189 177 0 3 22
0 21 27 25
0
0 0 624 0
6 74LS86
-21 -24 21 -16
3 U3C
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 3 0
1 U
3834 0 0
0
0
9 2-In XOR~
219 191 136 0 3 22
0 22 27 26
0
0 0 624 0
6 74LS86
-21 -24 21 -16
3 U3D
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 3 0
1 U
3363 0 0
0
0
6 74LS83
105 329 111 0 14 29
0 18 2 2 18 26 25 24 23 27
13 14 15 16 3
0
0 0 13040 0
7 74LS83A
-24 -60 25 -52
2 U4
-7 -61 7 -53
0
15 DVCC=5;DGND=12;
125 %D [%5bi %12bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 3 8 10 16 4 7 11 13
15 2 6 9 14 1 3 8 10 16
4 7 11 13 15 2 6 9 14 0
65 0 0 0 1 0 0 0
1 U
7668 0 0
0
0
9 V Source~
197 166 62 0 2 5
0 18 2
0
0 0 17264 0
3 10V
13 0 34 8
3 Vs1
13 -10 34 -2
0
0
11 %D %1 %2 %V
0
0
0
5

0 1 2 1 2 0
86 0 0 0 1 0 0 0
2 Vs
4718 0 0
0
0
7 Ground~
168 220 92 0 1 3
0 2
0
0 0 53360 0
0
4 GND5
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3874 0 0
0
0
9 Inverter~
13 417 61 0 2 22
0 13 10
0
0 0 624 0
6 74LS04
-21 -19 21 -11
2 s4
-8 -20 6 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 11 10 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 5 2 0
1 U
6671 0 0
0
0
9 Inverter~
13 419 98 0 2 22
0 14 9
0
0 0 624 0
6 74LS04
-21 -19 21 -11
2 s3
-8 -20 6 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 13 12 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 6 2 0
1 U
3789 0 0
0
0
9 Inverter~
13 421 139 0 2 22
0 15 8
0
0 0 624 0
6 74LS04
-21 -19 21 -11
2 s2
-10 -19 4 -11
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 4 0
1 U
4871 0 0
0
0
9 Inverter~
13 421 176 0 2 22
0 16 7
0
0 0 624 0
6 74LS04
-21 -19 21 -11
2 s1
-8 -20 6 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 4 0
1 U
3750 0 0
0
0
9 Inverter~
13 424 251 0 2 22
0 3 17
0
0 0 624 0
6 74LS04
-21 -19 21 -11
1 C
-4 -20 3 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 4 0
1 U
8778 0 0
0
0
7 Ground~
168 523 257 0 1 3
0 2
0
0 0 53360 0
0
4 GND4
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
538 0 0
0
0
7 Ground~
168 612 117 0 1 3
0 2
0
0 0 53360 0
0
4 GND6
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
6843 0 0
0
0
9 2-In AND~
219 636 187 0 3 22
0 4 3 6
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U6C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 5 0
1 U
3136 0 0
0
0
5 Lamp~
206 791 174 0 2 3
11 6 2
0
0 0 624 0
3 100
-10 -24 11 -16
1 Z
-4 -22 3 -14
0
0
11 %D %1 %2 %V
0
0
0
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 L
5950 0 0
0
0
5 Lamp~
206 515 238 0 2 3
11 17 2
0
0 0 624 0
3 100
-10 -24 11 -16
1 Y
-4 -20 3 -12
0
0
11 %D %1 %2 %V
0
0
0
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 L
5670 0 0
0
0
5 Lamp~
206 600 99 0 2 3
11 5 2
0
0 0 624 0
3 100
-10 -24 11 -16
1 X
-4 -21 3 -13
0
0
11 %D %1 %2 %V
0
0
0
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 L
6828 0 0
0
0
38
0 2 3 0 0 4224 0 0 25 19 0 2
369 196
612 196
2 1 4 0 0 8320 0 6 25 0 0 5
580 177
580 181
604 181
604 178
612 178
0 1 5 0 0 4224 0 0 6 12 0 2
580 112
580 141
3 1 6 0 0 4224 0 25 26 0 0 2
657 187
779 187
2 2 7 0 0 4224 0 21 7 0 0 4
442 176
465 176
465 164
473 164
2 1 8 0 0 4224 0 20 7 0 0 4
442 139
465 139
465 146
473 146
2 2 9 0 0 4224 0 19 8 0 0 4
440 98
462 98
462 87
470 87
2 1 10 0 0 4224 0 18 8 0 0 4
438 61
462 61
462 69
470 69
3 2 11 0 0 8320 0 7 9 0 0 6
518 155
522 155
522 131
518 131
518 121
523 121
3 1 12 0 0 8320 0 8 9 0 0 4
515 78
519 78
519 103
523 103
1 2 2 0 0 4096 0 10 26 0 0 2
803 191
803 187
3 1 5 0 0 0 0 9 28 0 0 4
568 112
566 112
566 112
588 112
1 2 2 0 0 0 0 24 28 0 0 2
612 111
612 112
10 1 13 0 0 8320 0 15 18 0 0 4
361 102
385 102
385 61
402 61
11 1 14 0 0 4224 0 15 19 0 0 4
361 111
396 111
396 98
404 98
12 1 15 0 0 4224 0 15 20 0 0 4
361 120
398 120
398 139
406 139
13 1 16 0 0 8320 0 15 21 0 0 4
361 129
385 129
385 176
406 176
2 1 17 0 0 4224 0 22 27 0 0 2
445 251
503 251
14 1 3 0 0 128 0 15 22 0 0 4
361 156
369 156
369 251
409 251
1 2 2 0 0 0 0 23 27 0 0 2
523 251
527 251
0 3 2 0 0 8192 0 0 15 22 0 3
270 84
270 93
297 93
0 2 2 0 0 8320 0 0 15 38 0 3
218 81
218 84
297 84
0 4 18 0 0 4096 0 0 15 24 0 3
257 37
257 102
297 102
1 1 18 0 0 8320 0 16 15 0 0 5
166 41
166 37
289 37
289 75
297 75
1 1 19 0 0 8320 0 2 11 0 0 5
84 294
84 253
162 253
162 254
170 254
1 1 20 0 0 8320 0 3 12 0 0 5
82 244
82 213
165 213
165 212
173 212
1 1 21 0 0 8320 0 4 13 0 0 3
79 186
79 168
173 168
1 1 22 0 0 4224 0 5 14 0 0 4
78 129
167 129
167 127
175 127
8 3 23 0 0 8320 0 15 11 0 0 4
297 138
266 138
266 263
219 263
7 3 24 0 0 8320 0 15 12 0 0 4
297 129
247 129
247 221
222 221
3 6 25 0 0 12416 0 13 15 0 0 4
222 177
236 177
236 120
297 120
3 5 26 0 0 8320 0 14 15 0 0 3
224 136
224 111
297 111
2 0 27 0 0 4096 0 11 0 0 36 2
170 272
116 272
2 0 27 0 0 4096 0 12 0 0 36 2
173 230
116 230
2 0 27 0 0 0 0 13 0 0 36 2
173 186
116 186
2 0 27 0 0 8320 0 14 0 0 37 3
175 145
116 145
116 336
1 9 27 0 0 0 0 1 15 0 0 4
101 336
289 336
289 156
297 156
2 1 2 0 0 0 0 16 17 0 0 6
166 83
166 88
207 88
207 81
220 81
220 86
4
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
521 222 553 246
531 230 555 246
3 A<B
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
798 161 830 185
808 169 832 185
3 A>B
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
609 82 641 106
619 90 643 106
3 A=B
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 4
109 47 149 71
119 55 151 71
4 1001
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
