CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 1 100 9
3 81 620 639
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
16 C:\CM60S\BOM.DAT
0 7
3 81 620 639
143654930 0
0
6 Title:
5 Name:
0
0
0
13
7 Ground~
168 469 94 0 1 3
0 2
0
0 0 53344 0
0
4 GND4
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
8953 0 0
0
0
7 Ground~
168 419 94 0 1 3
0 2
0
0 0 53344 0
0
4 GND3
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
4441 0 0
0
0
7 Ground~
168 359 97 0 1 3
0 2
0
0 0 53344 0
0
4 GND2
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3618 0 0
0
0
7 Ground~
168 302 96 0 1 3
0 2
0
0 0 53344 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
6153 0 0
0
0
6 74LS76
104 237 297 0 14 29
0 11 11 12 11 11 11 11 9 11
11 9 6 8 5
0
0 0 13024 0
6 74LS76
-21 -60 21 -52
2 U4
-7 -61 7 -53
0
15 DVCC=16;DGND=8;
131 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 4 16 1 2 3 9 12 6 7
8 15 14 11 10 4 16 1 2 3
9 12 6 7 8 15 14 11 10 0
65 0 0 0 1 0 0 0
1 U
5394 0 0
0
0
6 74LS76
104 411 297 0 14 29
0 10 10 8 10 10 10 10 7 10
10 7 4 13 3
0
0 0 13024 0
6 74LS76
-21 -60 21 -52
2 U5
-7 -61 7 -53
0
15 DVCC=16;DGND=8;
131 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 4 16 1 2 3 9 12 6 7
8 15 14 11 10 4 16 1 2 3
9 12 6 7 8 15 14 11 10 0
65 0 0 512 1 0 0 0
1 U
7734 0 0
0
0
7 Pulser~
4 61 352 0 10 12
0 14 15 12 16 0 0 5 5 1
7
0
0 0 4640 0
0
3 CLK
-10 -28 11 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
1 V
9914 0 0
0
0
2 +V
167 193 221 0 1 3
0 11
0
0 0 54240 0
2 5V
-7 -22 7 -14
2 V1
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
3747 0 0
0
0
2 +V
167 369 221 0 1 3
0 10
0
0 0 54240 0
2 5V
-7 -22 7 -14
2 V2
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
3549 0 0
0
0
5 Lamp~
206 459 75 0 2 3
11 6 2
0
0 0 624 0
3 100
-10 -24 11 -16
1 A
-4 -22 3 -14
0
0
11 %D %1 %2 %V
0
0
0
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 L
7931 0 0
0
0
5 Lamp~
206 406 75 0 2 3
11 5 2
0
0 0 624 0
3 100
-10 -24 11 -16
1 B
-4 -22 3 -14
0
0
11 %D %1 %2 %V
0
0
0
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 L
9325 0 0
0
0
5 Lamp~
206 347 77 0 2 3
11 4 2
0
0 0 624 0
3 100
-10 -24 11 -16
1 C
-4 -22 3 -14
0
0
11 %D %1 %2 %V
0
0
0
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 L
8903 0 0
0
0
5 Lamp~
206 291 77 0 2 3
11 3 2
0
0 0 624 0
3 100
-10 -24 11 -16
1 D
-4 -22 3 -14
0
0
11 %D %1 %2 %V
0
0
0
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 L
3834 0 0
0
0
28
1 2 2 0 0 4224 0 1 10 0 0 2
469 88
471 88
1 2 2 0 0 0 0 2 11 0 0 2
419 88
418 88
1 2 2 0 0 0 0 3 12 0 0 2
359 91
359 90
1 2 2 0 0 0 0 4 13 0 0 2
302 90
303 90
1 14 3 0 0 12416 0 13 6 0 0 6
279 90
275 90
275 114
489 114
489 315
449 315
12 1 4 0 0 8320 0 6 12 0 0 6
449 270
459 270
459 126
327 126
327 90
335 90
1 14 5 0 0 12416 0 11 5 0 0 5
394 88
394 158
309 158
309 315
275 315
12 1 6 0 0 12416 0 5 10 0 0 6
275 270
296 270
296 140
445 140
445 88
447 88
11 8 7 0 0 12416 0 6 6 0 0 6
443 261
468 261
468 366
347 366
347 324
373 324
13 3 8 0 0 4224 0 5 6 0 0 4
269 306
346 306
346 279
373 279
11 8 9 0 0 12416 0 5 5 0 0 6
269 261
287 261
287 367
178 367
178 324
199 324
1 0 10 0 0 4096 0 6 0 0 19 2
379 261
369 261
2 0 10 0 0 0 0 6 0 0 19 2
379 270
369 270
4 0 10 0 0 0 0 6 0 0 19 2
373 288
369 288
5 0 10 0 0 0 0 6 0 0 19 2
373 297
369 297
9 0 10 0 0 0 0 6 0 0 17 2
373 333
369 333
10 0 10 0 0 8192 0 6 0 0 19 3
373 342
369 342
369 315
6 0 10 0 0 0 0 6 0 0 19 2
379 306
369 306
7 1 10 0 0 8320 0 6 9 0 0 3
379 315
369 315
369 230
1 0 11 0 0 4096 0 5 0 0 27 2
205 261
193 261
2 0 11 0 0 0 0 5 0 0 27 2
205 270
193 270
4 0 11 0 0 0 0 5 0 0 27 2
199 288
193 288
5 0 11 0 0 0 0 5 0 0 27 2
199 297
193 297
9 0 11 0 0 0 0 5 0 0 25 2
199 333
193 333
10 0 11 0 0 8192 0 5 0 0 27 3
199 342
193 342
193 315
6 0 11 0 0 0 0 5 0 0 27 2
205 306
193 306
7 1 11 0 0 8320 0 5 8 0 0 3
205 315
193 315
193 230
3 3 12 0 0 12416 0 7 5 0 0 4
85 343
117 343
117 279
199 279
0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 100 100 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
12385 0
0 0.05 2
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
