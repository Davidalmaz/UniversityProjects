CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 9
32 88 1248 655
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
16 C:\CM60S\BOM.DAT
0 7
32 88 1248 655
143654930 0
0
6 Title:
5 Name:
0
0
0
11
13 Logic Switch~
5 278 321 0 10 11
0 7 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
1 D
-3 -26 4 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
8953 0 0
0
0
13 Logic Switch~
5 277 269 0 10 11
0 9 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
1 C
-3 -26 4 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
4441 0 0
0
0
13 Logic Switch~
5 278 210 0 1 11
0 8
0
0 0 21360 0
2 0V
-6 -16 8 -8
1 B
-3 -26 4 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
3618 0 0
0
0
13 Logic Switch~
5 280 137 0 1 11
0 11
0
0 0 21360 0
2 0V
-6 -16 8 -8
1 A
-3 -26 4 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
6153 0 0
0
0
7 Ground~
168 627 255 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
5394 0 0
0
0
10 3-In NAND~
219 578 249 0 4 22
0 6 4 5 3
0
0 0 624 0
6 74LS10
-21 -28 21 -20
3 U2A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
17

0 1 2 13 12 1 2 13 12 3
4 5 6 9 10 11 8 0
65 0 0 0 3 1 2 0
1 U
7734 0 0
0
0
10 2-In NAND~
219 451 312 0 3 22
0 8 7 5
0
0 0 624 0
6 74LS00
-14 -24 28 -16
3 U1D
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 1 0
1 U
9914 0 0
0
0
10 2-In NAND~
219 454 248 0 3 22
0 8 9 4
0
0 0 624 0
6 74LS00
-14 -24 28 -16
3 U1C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 1 0
1 U
3747 0 0
0
0
10 2-In NAND~
219 451 147 0 3 22
0 11 10 6
0
0 0 624 0
6 74LS00
-14 -24 28 -16
3 U1B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 1 0
1 U
3549 0 0
0
0
10 2-In NAND~
219 355 207 0 3 22
0 8 8 10
0
0 0 624 0
6 74LS00
-14 -24 28 -16
3 U1A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 1 0
1 U
7931 0 0
0
0
5 Lamp~
206 615 236 0 2 3
11 3 2
0
0 0 608 0
3 100
-10 -24 11 -16
2 L1
-7 -22 7 -14
0
0
11 %D %1 %2 %V
0
0
0
5

0 1 2 1 2 0
82 0 0 0 0 0 0 0
1 L
9325 0 0
0
0
13
1 2 2 0 0 0 0 5 11 0 0 2
627 249
627 249
1 4 3 0 0 4224 0 11 6 0 0 2
603 249
605 249
3 2 4 0 0 4224 0 8 6 0 0 4
481 248
544 248
544 249
554 249
3 3 5 0 0 4224 0 7 6 0 0 4
478 312
544 312
544 258
554 258
3 1 6 0 0 8320 0 9 6 0 0 4
478 147
544 147
544 240
554 240
1 2 7 0 0 4224 0 1 7 0 0 2
290 321
427 321
0 1 8 0 0 8320 0 0 7 12 0 3
298 210
298 303
427 303
1 2 9 0 0 4224 0 2 8 0 0 4
289 269
422 269
422 257
430 257
0 1 8 0 0 0 0 0 8 12 0 3
313 210
313 239
430 239
3 2 10 0 0 8320 0 10 9 0 0 4
382 207
419 207
419 156
427 156
0 2 8 0 0 0 0 0 10 12 0 3
323 210
323 216
331 216
1 1 8 0 0 0 0 3 10 0 0 4
290 210
323 210
323 198
331 198
1 1 11 0 0 4224 0 4 9 0 0 4
292 137
418 137
418 138
427 138
0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
