CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 80 9
0 71 1280 672
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
16 C:\CM60S\BOM.DAT
0 7
0 71 1280 672
143654930 0
0
6 Title:
5 Name:
0
0
0
44
7 Ground~
168 394 26 0 1 3
0 0
0
0 0 53344 180
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
8953 0 0
0
0
13 Logic Switch~
5 22 328 0 10 11
0 2 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
3 V29
-9 -26 12 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
4441 0 0
0
0
13 Logic Switch~
5 23 290 0 10 11
0 3 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
3 V28
-9 -26 12 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
3618 0 0
0
0
13 Logic Switch~
5 26 207 0 1 11
0 5
0
0 0 21360 0
2 0V
-6 -16 8 -8
3 V27
-9 -26 12 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
6153 0 0
0
0
13 Logic Switch~
5 26 248 0 10 11
0 4 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
3 V26
-9 -26 12 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
5394 0 0
0
0
13 Logic Switch~
5 83 666 0 10 11
0 8 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
3 V25
-9 -26 12 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
7734 0 0
0
0
13 Logic Switch~
5 83 625 0 1 11
0 9
0
0 0 21360 0
2 0V
-6 -16 8 -8
3 V24
-9 -26 12 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
9914 0 0
0
0
13 Logic Switch~
5 80 708 0 10 11
0 7 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
3 V23
-9 -26 12 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
3747 0 0
0
0
13 Logic Switch~
5 79 746 0 1 11
0 6
0
0 0 21360 0
2 0V
-6 -16 8 -8
3 V17
-9 -26 12 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3549 0 0
0
0
13 Logic Switch~
5 83 568 0 10 11
0 10 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
3 V12
-9 -26 12 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
7931 0 0
0
0
13 Logic Switch~
5 84 530 0 1 11
0 11
0
0 0 21360 0
2 0V
-6 -16 8 -8
3 V11
-9 -26 12 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
9325 0 0
0
0
13 Logic Switch~
5 87 447 0 1 11
0 13
0
0 0 21360 0
2 0V
-6 -16 8 -8
3 V10
-9 -26 12 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
8903 0 0
0
0
13 Logic Switch~
5 87 488 0 10 11
0 12 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V9
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
3834 0 0
0
0
13 Logic Switch~
5 491 42 0 10 11
0 14 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
1 Z
-3 -26 4 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3363 0 0
0
0
13 Logic Switch~
5 90 307 0 10 11
0 17 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V8
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
7668 0 0
0
0
13 Logic Switch~
5 90 266 0 1 11
0 18
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V7
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
4718 0 0
0
0
13 Logic Switch~
5 87 349 0 1 11
0 16
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V6
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3874 0 0
0
0
13 Logic Switch~
5 86 387 0 1 11
0 15
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V5
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
6671 0 0
0
0
13 Logic Switch~
5 601 523 0 1 11
0 30
0
0 0 21360 0
2 0V
-6 -16 8 -8
3 V15
-9 -26 12 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3789 0 0
0
0
13 Logic Switch~
5 604 440 0 1 11
0 28
0
0 0 21360 0
2 0V
-6 -16 8 -8
3 V14
-9 -26 12 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
4871 0 0
0
0
13 Logic Switch~
5 604 481 0 1 11
0 29
0
0 0 21360 0
2 0V
-6 -16 8 -8
3 V13
-9 -26 12 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3750 0 0
0
0
13 Logic Switch~
5 389 319 0 1 11
0 34
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V4
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
8778 0 0
0
0
13 Logic Switch~
5 389 278 0 1 11
0 35
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V3
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
538 0 0
0
0
13 Logic Switch~
5 384 365 0 10 11
0 33 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
6843 0 0
0
0
13 Logic Switch~
5 383 403 0 1 11
0 32
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3136 0 0
0
0
13 Logic Switch~
5 817 737 0 1 11
0 27
0
0 0 21360 0
2 0V
-6 -16 8 -8
3 V33
-9 -26 12 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5950 0 0
0
0
13 Logic Switch~
5 818 699 0 1 11
0 26
0
0 0 21360 0
2 0V
-6 -16 8 -8
3 V32
-9 -26 12 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5670 0 0
0
0
13 Logic Switch~
5 821 616 0 1 11
0 24
0
0 0 21360 0
2 0V
-6 -16 8 -8
3 V31
-9 -26 12 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
6828 0 0
0
0
13 Logic Switch~
5 821 657 0 1 11
0 25
0
0 0 21360 0
2 0V
-6 -16 8 -8
3 V30
-9 -26 12 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
6735 0 0
0
0
13 Logic Switch~
5 549 42 0 10 11
0 41 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
1 X
-3 -26 4 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
8365 0 0
0
0
13 Logic Switch~
5 647 48 0 10 11
0 40 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
1 W
-3 -26 4 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
4132 0 0
0
0
13 Logic Switch~
5 601 557 0 10 11
0 31 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
3 V16
-9 -26 12 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
4551 0 0
0
0
13 Logic Switch~
5 92 162 0 10 11
0 36 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
3 V19
-9 -26 12 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
3635 0 0
0
0
13 Logic Switch~
5 93 124 0 10 11
0 38 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
3 V20
-9 -26 12 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
3973 0 0
0
0
13 Logic Switch~
5 96 41 0 1 11
0 39
0
0 0 21360 0
2 0V
-6 -16 8 -8
3 V21
-9 -26 12 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3851 0 0
0
0
13 Logic Switch~
5 96 82 0 1 11
0 37
0
0 0 21360 0
2 0V
-6 -16 8 -8
3 V22
-9 -26 12 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
8383 0 0
0
0
7 74LS151
20 981 677 0 14 29
0 2 6 10 15 36 32 31 27 42
14 41 40 19 51
0
0 0 13040 0
7 74LS151
-24 -60 25 -52
7 William
-24 -61 25 -53
0
15 DVCC=16;DGND=8;
141 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i %12i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 12 13 14 15 1 2 3 4 7
9 10 11 5 6 12 13 14 15 1
2 3 4 7 9 10 11 5 6 0
65 0 0 512 1 0 0 0
1 U
9334 0 0
0
0
7 74LS151
20 704 490 0 14 29
0 3 7 11 16 38 33 30 26 42
14 41 40 20 52
0
0 0 13040 0
7 74LS151
-24 -60 25 -52
6 Xavier
-21 -61 21 -53
0
15 DVCC=16;DGND=8;
141 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i %12i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 12 13 14 15 1 2 3 4 7
9 10 11 5 6 12 13 14 15 1
2 3 4 7 9 10 11 5 6 0
65 0 0 512 1 0 0 0
1 U
7471 0 0
0
0
7 74LS151
20 497 336 0 14 29
0 4 8 12 17 37 34 29 25 42
14 41 40 21 53
0
0 0 13040 0
7 74LS151
-24 -60 25 -52
7 Yelitza
-24 -61 25 -53
0
15 DVCC=16;DGND=8;
141 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i %12i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 12 13 14 15 1 2 3 4 7
9 10 11 5 6 12 13 14 15 1
2 3 4 7 9 10 11 5 6 0
65 0 0 512 1 0 0 0
1 U
3334 0 0
0
0
2 +V
167 1307 87 0 1 3
0 50
0
0 0 54256 0
2 5V
-7 -22 7 -14
3 V18
-10 -32 11 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
3559 0 0
0
0
6 74LS47
187 1091 224 0 14 29
0 22 21 20 19 54 55 43 44 45
46 47 48 49 56
0
0 0 13040 0
6 74LS47
-21 -60 21 -52
2 U1
-7 -61 7 -53
0
15 DVCC=16;DGND=8;
119 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %14i]
+ [%16bo %1o %2o %3o %4o %5o %6o %14o %7o %8o %9o %10o %11o %12o %13o] %M
0
12 type:digital
5 DIP16
29

0 6 2 1 7 3 5 14 15 9
10 11 12 13 4 6 2 1 7 3
5 14 15 9 10 11 12 13 4 0
65 0 0 512 1 0 0 0
1 U
984 0 0
0
0
9 CA 7-Seg~
184 1215 149 0 18 19
10 49 48 47 46 45 44 43 57 23
0 0 0 2 2 2 2 2 1
0
0 0 21104 0
5 REDCA
16 -41 51 -33
5 DISP2
30 -4 65 4
0
0
32 %D %1 %2 %3 %4 %5 %6 %7 %8 %9 %S
0
0
0
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
88 0 0 512 1 0 0 0
4 DISP
7557 0 0
0
0
7 74LS151
20 326 103 0 14 29
0 5 9 13 18 39 35 28 24 42
14 41 40 22 58
0
0 0 13040 0
7 74LS151
-24 -60 25 -52
5 Zaida
-17 -61 18 -53
0
15 DVCC=16;DGND=8;
141 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i %12i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 12 13 14 15 1 2 3 4 7
9 10 11 5 6 12 13 14 15 1
2 3 4 7 9 10 11 5 6 0
65 0 0 512 1 0 0 0
1 U
3146 0 0
0
0
9 Resistor~
219 1263 99 0 4 5
0 23 50 0 1
0
0 0 880 0
6 0.047k
-20 -14 22 -6
2 R2
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
5687 0 0
0
0
61
1 1 2 0 0 12416 0 2 37 0 0 6
34 328
369 328
369 668
941 668
941 650
949 650
1 1 3 0 0 4224 0 3 38 0 0 4
35 290
461 290
461 463
672 463
1 1 4 0 0 4224 0 5 39 0 0 4
38 248
457 248
457 309
465 309
1 1 5 0 0 4224 0 4 43 0 0 4
38 207
286 207
286 76
294 76
1 2 6 0 0 4224 0 9 37 0 0 6
91 746
803 746
803 646
941 646
941 659
949 659
1 2 7 0 0 4224 0 8 38 0 0 4
92 708
664 708
664 472
672 472
1 2 8 0 0 4224 0 6 39 0 0 4
95 666
457 666
457 318
465 318
1 2 9 0 0 8320 0 7 43 0 0 4
95 625
286 625
286 85
294 85
1 3 10 0 0 4224 0 10 37 0 0 4
95 568
941 568
941 668
949 668
1 3 11 0 0 4224 0 11 38 0 0 6
96 530
587 530
587 470
664 470
664 481
672 481
1 3 12 0 0 4224 0 13 39 0 0 4
99 488
457 488
457 327
465 327
1 3 13 0 0 8320 0 12 43 0 0 4
99 447
286 447
286 94
294 94
0 1 14 0 0 4096 0 0 14 49 0 3
512 86
512 42
503 42
1 4 15 0 0 4224 0 18 37 0 0 4
98 387
941 387
941 677
949 677
1 4 16 0 0 4224 0 17 38 0 0 5
99 349
461 349
461 491
672 491
672 490
1 4 17 0 0 4240 0 15 39 0 0 4
102 307
457 307
457 336
465 336
1 4 18 0 0 4224 0 16 43 0 0 6
102 266
294 266
294 153
286 153
286 103
294 103
4 13 19 0 0 8320 0 41 37 0 0 4
1059 215
1027 215
1027 704
1013 704
3 13 20 0 0 8320 0 41 38 0 0 4
1059 206
750 206
750 517
736 517
2 13 21 0 0 4224 0 41 39 0 0 4
1059 197
543 197
543 363
529 363
1 13 22 0 0 4224 0 41 43 0 0 4
1059 188
372 188
372 130
358 130
1 9 23 0 0 4224 0 44 42 0 0 3
1245 99
1215 99
1215 113
1 8 24 0 0 12416 0 28 43 0 0 6
833 616
868 616
868 164
286 164
286 139
294 139
1 8 25 0 0 12416 0 29 39 0 0 6
833 657
850 657
850 387
457 387
457 372
465 372
1 8 26 0 0 12416 0 27 38 0 0 6
830 699
839 699
839 541
664 541
664 526
672 526
1 8 27 0 0 4224 0 26 37 0 0 5
829 737
941 737
941 712
949 712
949 713
1 7 28 0 0 12416 0 20 43 0 0 6
616 440
621 440
621 155
286 155
286 130
294 130
1 7 29 0 0 12416 0 21 39 0 0 6
616 481
621 481
621 387
457 387
457 363
465 363
1 7 30 0 0 4224 0 19 38 0 0 4
613 523
664 523
664 517
672 517
1 7 31 0 0 4224 0 32 37 0 0 5
613 557
931 557
931 703
949 703
949 704
1 6 32 0 0 4224 0 25 37 0 0 5
395 403
875 403
875 694
949 694
949 695
1 6 33 0 0 12416 0 24 38 0 0 4
396 365
461 365
461 508
672 508
1 6 34 0 0 4224 0 22 39 0 0 4
401 319
457 319
457 354
465 354
1 6 35 0 0 12416 0 23 43 0 0 6
401 278
406 278
406 170
262 170
262 121
294 121
1 5 36 0 0 12416 0 33 37 0 0 5
104 162
134 162
134 685
949 685
949 686
1 5 37 0 0 8320 0 36 39 0 0 4
108 82
226 82
226 345
465 345
1 5 38 0 0 12416 0 34 38 0 0 4
105 124
184 124
184 499
672 499
1 5 39 0 0 4224 0 35 43 0 0 4
108 41
258 41
258 112
294 112
12 0 40 0 0 16512 0 37 0 0 44 5
1013 677
1013 676
1306 676
1306 604
983 604
11 0 41 0 0 16512 0 37 0 0 45 5
1013 668
1013 667
1286 667
1286 570
957 570
10 0 14 0 0 16512 0 37 0 0 46 5
1013 659
1013 658
1254 658
1254 556
939 556
9 0 42 0 0 16512 0 37 0 0 43 5
1019 650
1019 649
1230 649
1230 546
913 546
9 0 42 0 0 0 0 38 0 0 50 6
742 463
913 463
913 546
913 546
913 300
642 300
12 0 40 0 0 0 0 38 0 0 47 6
736 490
983 490
983 604
983 604
983 351
771 351
11 0 41 0 0 0 0 38 0 0 48 6
736 481
957 481
957 570
957 570
957 331
735 331
10 0 14 0 0 0 0 38 0 0 49 6
736 472
939 472
939 556
939 556
939 321
700 321
12 0 40 0 0 0 0 39 0 0 51 6
529 336
771 336
771 351
771 351
771 75
668 75
11 0 41 0 0 0 0 39 0 0 52 6
529 327
735 327
735 335
735 335
735 62
570 62
10 10 14 0 0 0 0 39 43 0 0 6
529 318
700 318
700 86
490 86
490 85
358 85
9 0 42 0 0 0 0 39 0 0 53 4
535 309
642 309
642 76
395 76
12 1 40 0 0 0 0 43 31 0 0 4
358 103
668 103
668 48
659 48
11 1 41 0 0 0 0 43 30 0 0 4
358 94
570 94
570 42
561 42
9 1 42 0 0 0 0 43 1 0 0 4
364 76
395 76
395 34
394 34
7 7 43 0 0 8320 0 42 41 0 0 3
1230 185
1230 188
1129 188
6 8 44 0 0 8320 0 42 41 0 0 3
1224 185
1224 197
1129 197
5 9 45 0 0 8320 0 42 41 0 0 3
1218 185
1218 206
1129 206
4 10 46 0 0 8320 0 42 41 0 0 3
1212 185
1212 215
1129 215
3 11 47 0 0 8320 0 42 41 0 0 3
1206 185
1206 224
1129 224
2 12 48 0 0 8320 0 42 41 0 0 3
1200 185
1200 233
1129 233
1 13 49 0 0 8320 0 42 41 0 0 3
1194 185
1194 242
1129 242
2 1 50 0 0 4224 0 44 40 0 0 3
1281 99
1307 99
1307 96
0
0
2065 0 1
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 5e-006 2e-008 2e-008
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
1181856 1079360 100 100 0 0
0 0 0 0
0 71 161 141
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
12385 0
4 1 2
0
9634944 8550464 100 100 0 0
77 66 1247 216
0 371 1280 671
1247 66
77 66
1247 66
1247 216
0 0
0 0 0 0 0 0
12385 0
4 1e-006 2
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
