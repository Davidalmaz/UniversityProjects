CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 5 100 9
38 96 1498 799
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
16 C:\CM60S\BOM.DAT
0 7
38 588 1498 799
160432146 0
0
6 Title:
5 Name:
0
0
0
9
5 SCOPE
12 562 335 0 1 11
0 2
0
0 0 57568 0
3 SAL
-11 -4 10 4
2 U1
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
0
8953 0 0
0
0
5 SCOPE
12 195 113 0 1 11
0 2
0
0 0 57584 0
3 ENT
-11 -4 10 4
2 U1
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
0
4441 0 0
0
0
7 Pulser~
4 135 133 0 10 12
0 9 10 2 11 0 0 5 5 1
8
0
0 0 4656 0
0
5 PULSO
-17 -28 18 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 0 0 0 0
1 V
3618 0 0
0
0
9 Inverter~
13 518 346 0 2 22
0 4 3
0
0 0 624 0
6 74LS04
-21 -19 21 -11
4 NOT6
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
15

0 13 12 1 2 3 4 5 6 9
8 11 10 13 12 0
65 0 0 0 6 6 1 0
1 U
6153 0 0
0
0
9 Inverter~
13 460 304 0 2 22
0 5 4
0
0 0 624 0
6 74LS04
-21 -19 21 -11
4 NOT5
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
15

0 11 10 1 2 3 4 5 6 9
8 11 10 13 12 0
65 0 0 0 6 5 1 0
1 U
5394 0 0
0
0
9 Inverter~
13 398 258 0 2 22
0 6 5
0
0 0 624 0
6 74LS04
-21 -19 21 -11
4 NOT4
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
15

0 9 8 1 2 3 4 5 6 9
8 11 10 13 12 0
65 0 0 0 6 4 1 0
1 U
7734 0 0
0
0
9 Inverter~
13 346 215 0 2 22
0 7 6
0
0 0 624 0
6 74LS04
-21 -19 21 -11
4 NOT3
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
15

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0
65 0 0 0 6 3 1 0
1 U
9914 0 0
0
0
9 Inverter~
13 292 173 0 2 22
0 8 7
0
0 0 624 0
6 74LS04
-21 -19 21 -11
4 NOT2
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
15

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0
65 0 0 0 6 2 1 0
1 U
3747 0 0
0
0
9 Inverter~
13 242 125 0 2 22
0 2 8
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 NOT
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
15

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0
65 0 0 0 6 1 1 0
1 U
3549 0 0
0
0
8
1 0 2 0 0 0 0 2 0 0 3 2
195 125
195 125
2 1 3 0 0 4224 0 4 1 0 0 3
539 346
562 346
562 347
3 1 2 0 0 4224 0 3 9 0 0 4
159 124
195 124
195 125
227 125
2 1 4 0 0 8320 0 5 4 0 0 4
481 304
502 304
502 346
503 346
2 1 5 0 0 8320 0 6 5 0 0 4
419 258
437 258
437 304
445 304
2 1 6 0 0 8320 0 7 6 0 0 4
367 215
375 215
375 258
383 258
2 1 7 0 0 8320 0 8 7 0 0 4
313 173
323 173
323 215
331 215
2 1 8 0 0 8320 0 9 8 0 0 4
263 125
269 125
269 173
277 173
0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 100 100 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
12385 0
0 2 2
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
