CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 5 100 9
14 83 687 795
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
16 C:\CM60S\BOM.DAT
0 7
35 606 708 747
160432146 0
0
6 Title:
5 Name:
0
0
0
8
9 2-In XOR~
219 456 106 0 3 22
0 6 4 3
0
0 0 624 0
6 74LS86
-21 -24 21 -16
3 U1A
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 1 0
1 U
8953 0 0
0
0
5 SCOPE
12 520 94 0 1 11
0 3
0
0 0 57584 0
3 SAL
-11 -4 10 4
2 U2
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
0
4441 0 0
0
0
5 SCOPE
12 364 121 0 1 11
0 4
0
0 0 57584 0
2 E1
-7 -4 7 4
2 U2
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
0
3618 0 0
0
0
5 SCOPE
12 364 95 0 1 11
0 6
0
0 0 57584 0
2 E2
-8 -4 6 4
2 U2
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
0
6153 0 0
0
0
7 Ground~
168 337 181 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
5394 0 0
0
0
7 Pulser~
4 100 115 0 10 12
0 7 8 5 9 0 0 5 5 4
7
0
0 0 4656 0
0
5 RELOJ
-17 -28 18 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
1 V
7734 0 0
0
0
6 74LS93
109 256 97 0 8 17
0 2 2 5 4 10 11 6 4
0
0 0 13040 0
6 74LS93
-21 -35 21 -27
4 CONT
-14 -36 14 -28
0
15 DVCC=5;DGND=10;
76 %D [%5bi %10bi %1i %2i %3i %4i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o] %M
0
12 type:digital
5 DIP14
17

0 2 3 14 1 11 8 9 12 2
3 14 1 11 8 9 12 0
65 0 0 512 1 0 0 0
1 U
9914 0 0
0
0
5 Lamp~
206 570 92 0 2 3
11 3 2
0
0 0 608 0
3 100
-10 -24 11 -16
4 LAMP
-14 -22 14 -14
0
0
11 %D %1 %2 %V
0
0
0
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 L
3747 0 0
0
0
12
2 1 2 0 0 12416 0 8 5 0 0 5
582 105
586 105
586 167
337 167
337 175
3 0 3 0 0 4096 0 1 0 0 12 2
489 106
489 105
4 8 4 0 0 12288 0 7 7 0 0 5
218 115
214 115
214 144
288 144
288 115
3 3 5 0 0 4224 0 6 7 0 0 2
124 106
218 106
1 0 3 0 0 0 0 2 0 0 12 2
520 106
520 105
1 0 4 0 0 0 0 3 0 0 9 2
364 133
364 134
1 0 6 0 0 4096 0 4 0 0 8 2
364 107
364 106
7 1 6 0 0 4224 0 7 1 0 0 7
288 106
431 106
431 96
438 96
438 96
440 96
440 97
8 2 4 0 0 12416 0 7 1 0 0 9
288 115
300 115
300 134
431 134
431 114
438 114
438 114
440 114
440 115
2 0 2 0 0 0 0 7 0 0 11 2
224 97
200 97
1 1 2 0 0 0 0 7 5 0 0 5
224 88
200 88
200 167
337 167
337 175
0 1 3 0 0 4224 0 0 8 0 0 2
482 105
558 105
0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
