CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 5 100 9
0 71 1280 680
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
16 C:\CM60S\BOM.DAT
0 7
0 71 1280 680
143654930 0
0
6 Title:
5 Name:
0
0
0
10
13 Logic Switch~
5 251 219 0 10 11
0 6 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-7 -15 7 -7
1 C
-3 -26 4 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
8953 0 0
0
0
13 Logic Switch~
5 258 285 0 10 11
0 7 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-7 -15 7 -7
1 D
-3 -26 4 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
4441 0 0
0
0
13 Logic Switch~
5 252 133 0 10 11
0 8 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-7 -15 7 -7
1 B
-3 -26 4 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
3618 0 0
0
0
13 Logic Switch~
5 245 67 0 10 11
0 9 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-10 -14 4 -6
1 A
-3 -26 4 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
6153 0 0
0
0
7 Ground~
168 592 131 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
5394 0 0
0
0
10 2-In NAND~
219 463 185 0 3 22
0 10 11 12
0
0 0 112 0
6 74LS00
-14 -24 28 -16
0
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 512 4 1 2 0
1 U
7734 0 0
0
0
10 2-In NAND~
219 371 190 0 3 22
0 6 7 4
0
0 0 624 0
6 74LS00
-14 -24 28 -16
3 CDN
-4 -34 17 -26
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 2 0
1 U
9914 0 0
0
0
10 2-In NAND~
219 455 126 0 3 22
0 5 4 3
0
0 0 112 0
6 74LS00
-14 -24 28 -16
0
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 2 0
1 U
3747 0 0
0
0
10 2-In NAND~
219 375 123 0 3 22
0 9 8 5
0
0 0 624 0
6 74LS00
-14 -24 28 -16
3 ABN
-4 -34 17 -26
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 2 0
1 U
3549 0 0
0
0
5 Lamp~
206 580 112 0 2 3
11 3 2
0
0 0 624 0
3 100
-10 -24 11 -16
2 L1
-7 -22 7 -14
0
0
11 %D %1 %2 %V
0
0
0
5

0 1 2 1 2 0
82 0 0 0 0 0 0 0
1 L
7931 0 0
0
0
8
3 1 3 0 0 8320 0 8 10 0 0 3
482 126
482 125
568 125
3 2 4 0 0 8320 0 7 8 0 0 4
398 190
421 190
421 135
431 135
3 1 5 0 0 4224 0 9 8 0 0 4
402 123
423 123
423 117
431 117
1 1 6 0 0 8320 0 1 7 0 0 3
263 219
263 181
347 181
1 2 7 0 0 8320 0 2 7 0 0 4
270 285
339 285
339 199
347 199
1 2 8 0 0 4224 0 3 9 0 0 4
264 133
343 133
343 132
351 132
1 1 9 0 0 4224 0 4 9 0 0 4
257 67
343 67
343 114
351 114
1 2 2 0 0 0 0 5 10 0 0 2
592 125
592 125
1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 10
418 87 506 111
428 95 508 111
10 (Ab'*Cd')'
0
2049 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
788264 1079360 100 100 0 0
0 0 0 0
1 66 162 136
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
12385 0
4 2 2
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
